module tt_um_piggy_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire net32;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire net31;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire net30;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire net29;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire net28;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire clknet_leaf_0_clk;
 wire \ascii0[0] ;
 wire \ascii0[10] ;
 wire \ascii0[11] ;
 wire \ascii0[12] ;
 wire \ascii0[16] ;
 wire \ascii0[17] ;
 wire \ascii0[1] ;
 wire \ascii0[20] ;
 wire \ascii0[2] ;
 wire \ascii0[3] ;
 wire \ascii0[8] ;
 wire \ascii0[9] ;
 wire \ascii1[0] ;
 wire \ascii1[10] ;
 wire \ascii1[11] ;
 wire \ascii1[12] ;
 wire \ascii1[16] ;
 wire \ascii1[17] ;
 wire \ascii1[1] ;
 wire \ascii1[20] ;
 wire \ascii1[2] ;
 wire \ascii1[3] ;
 wire \ascii1[8] ;
 wire \ascii1[9] ;
 wire \ascii2[0] ;
 wire \ascii2[10] ;
 wire \ascii2[11] ;
 wire \ascii2[12] ;
 wire \ascii2[16] ;
 wire \ascii2[17] ;
 wire \ascii2[1] ;
 wire \ascii2[20] ;
 wire \ascii2[2] ;
 wire \ascii2[3] ;
 wire \ascii2[8] ;
 wire \ascii2[9] ;
 wire \ascii3[0] ;
 wire \ascii3[10] ;
 wire \ascii3[11] ;
 wire \ascii3[12] ;
 wire \ascii3[16] ;
 wire \ascii3[17] ;
 wire \ascii3[1] ;
 wire \ascii3[20] ;
 wire \ascii3[2] ;
 wire \ascii3[3] ;
 wire \ascii3[8] ;
 wire \ascii3[9] ;
 wire change0;
 wire change1;
 wire change2;
 wire change3;
 wire o_Tx_Active;
 wire o_Tx_Done;
 wire o_Tx_Serial;
 wire or4_out;
 wire start_sending;
 wire \u_cnt0.count[0] ;
 wire \u_cnt0.count[1] ;
 wire \u_cnt0.count[2] ;
 wire \u_cnt0.count[3] ;
 wire \u_cnt0.count[4] ;
 wire \u_cnt0.count[5] ;
 wire \u_cnt0.count[6] ;
 wire \u_cnt0.count[7] ;
 wire \u_cnt0.state ;
 wire \u_cnt1.count[0] ;
 wire \u_cnt1.count[1] ;
 wire \u_cnt1.count[2] ;
 wire \u_cnt1.count[3] ;
 wire \u_cnt1.count[4] ;
 wire \u_cnt1.count[5] ;
 wire \u_cnt1.count[6] ;
 wire \u_cnt1.count[7] ;
 wire \u_cnt1.state ;
 wire \u_cnt2.count[0] ;
 wire \u_cnt2.count[1] ;
 wire \u_cnt2.count[2] ;
 wire \u_cnt2.count[3] ;
 wire \u_cnt2.count[4] ;
 wire \u_cnt2.count[5] ;
 wire \u_cnt2.count[6] ;
 wire \u_cnt2.count[7] ;
 wire \u_cnt2.state ;
 wire \u_cnt3.count[0] ;
 wire \u_cnt3.count[1] ;
 wire \u_cnt3.count[2] ;
 wire \u_cnt3.count[3] ;
 wire \u_cnt3.count[4] ;
 wire \u_cnt3.count[5] ;
 wire \u_cnt3.count[6] ;
 wire \u_cnt3.count[7] ;
 wire \u_cnt3.state ;
 wire \u_deb0.Output ;
 wire \u_deb0.counter[0] ;
 wire \u_deb0.counter[10] ;
 wire \u_deb0.counter[11] ;
 wire \u_deb0.counter[12] ;
 wire \u_deb0.counter[13] ;
 wire \u_deb0.counter[14] ;
 wire \u_deb0.counter[15] ;
 wire \u_deb0.counter[16] ;
 wire \u_deb0.counter[17] ;
 wire \u_deb0.counter[18] ;
 wire \u_deb0.counter[19] ;
 wire \u_deb0.counter[1] ;
 wire \u_deb0.counter[2] ;
 wire \u_deb0.counter[3] ;
 wire \u_deb0.counter[4] ;
 wire \u_deb0.counter[5] ;
 wire \u_deb0.counter[6] ;
 wire \u_deb0.counter[7] ;
 wire \u_deb0.counter[8] ;
 wire \u_deb0.counter[9] ;
 wire \u_deb1.Output ;
 wire \u_deb1.counter[0] ;
 wire \u_deb1.counter[10] ;
 wire \u_deb1.counter[11] ;
 wire \u_deb1.counter[12] ;
 wire \u_deb1.counter[13] ;
 wire \u_deb1.counter[14] ;
 wire \u_deb1.counter[15] ;
 wire \u_deb1.counter[16] ;
 wire \u_deb1.counter[17] ;
 wire \u_deb1.counter[18] ;
 wire \u_deb1.counter[19] ;
 wire \u_deb1.counter[1] ;
 wire \u_deb1.counter[2] ;
 wire \u_deb1.counter[3] ;
 wire \u_deb1.counter[4] ;
 wire \u_deb1.counter[5] ;
 wire \u_deb1.counter[6] ;
 wire \u_deb1.counter[7] ;
 wire \u_deb1.counter[8] ;
 wire \u_deb1.counter[9] ;
 wire \u_deb2.Output ;
 wire \u_deb2.counter[0] ;
 wire \u_deb2.counter[10] ;
 wire \u_deb2.counter[11] ;
 wire \u_deb2.counter[12] ;
 wire \u_deb2.counter[13] ;
 wire \u_deb2.counter[14] ;
 wire \u_deb2.counter[15] ;
 wire \u_deb2.counter[16] ;
 wire \u_deb2.counter[17] ;
 wire \u_deb2.counter[18] ;
 wire \u_deb2.counter[19] ;
 wire \u_deb2.counter[1] ;
 wire \u_deb2.counter[2] ;
 wire \u_deb2.counter[3] ;
 wire \u_deb2.counter[4] ;
 wire \u_deb2.counter[5] ;
 wire \u_deb2.counter[6] ;
 wire \u_deb2.counter[7] ;
 wire \u_deb2.counter[8] ;
 wire \u_deb2.counter[9] ;
 wire \u_deb3.Output ;
 wire \u_deb3.counter[0] ;
 wire \u_deb3.counter[10] ;
 wire \u_deb3.counter[11] ;
 wire \u_deb3.counter[12] ;
 wire \u_deb3.counter[13] ;
 wire \u_deb3.counter[14] ;
 wire \u_deb3.counter[15] ;
 wire \u_deb3.counter[16] ;
 wire \u_deb3.counter[17] ;
 wire \u_deb3.counter[18] ;
 wire \u_deb3.counter[19] ;
 wire \u_deb3.counter[1] ;
 wire \u_deb3.counter[2] ;
 wire \u_deb3.counter[3] ;
 wire \u_deb3.counter[4] ;
 wire \u_deb3.counter[5] ;
 wire \u_deb3.counter[6] ;
 wire \u_deb3.counter[7] ;
 wire \u_deb3.counter[8] ;
 wire \u_deb3.counter[9] ;
 wire \u_deb4.Output ;
 wire \u_deb4.counter[0] ;
 wire \u_deb4.counter[10] ;
 wire \u_deb4.counter[11] ;
 wire \u_deb4.counter[12] ;
 wire \u_deb4.counter[13] ;
 wire \u_deb4.counter[14] ;
 wire \u_deb4.counter[15] ;
 wire \u_deb4.counter[16] ;
 wire \u_deb4.counter[17] ;
 wire \u_deb4.counter[18] ;
 wire \u_deb4.counter[19] ;
 wire \u_deb4.counter[1] ;
 wire \u_deb4.counter[2] ;
 wire \u_deb4.counter[3] ;
 wire \u_deb4.counter[4] ;
 wire \u_deb4.counter[5] ;
 wire \u_deb4.counter[6] ;
 wire \u_deb4.counter[7] ;
 wire \u_deb4.counter[8] ;
 wire \u_deb4.counter[9] ;
 wire \u_edge.Output ;
 wire \u_edge.state ;
 wire \u_n2a0.hundreds[0] ;
 wire \u_n2a0.hundreds[1] ;
 wire \u_n2a0.ones[0] ;
 wire \u_n2a0.ones[1] ;
 wire \u_n2a0.ones[2] ;
 wire \u_n2a0.ones[3] ;
 wire \u_n2a0.tens[0] ;
 wire \u_n2a0.tens[1] ;
 wire \u_n2a0.tens[2] ;
 wire \u_n2a0.tens[3] ;
 wire \u_n2a1.hundreds[0] ;
 wire \u_n2a1.hundreds[1] ;
 wire \u_n2a1.ones[0] ;
 wire \u_n2a1.ones[1] ;
 wire \u_n2a1.ones[2] ;
 wire \u_n2a1.ones[3] ;
 wire \u_n2a1.tens[0] ;
 wire \u_n2a1.tens[1] ;
 wire \u_n2a1.tens[2] ;
 wire \u_n2a1.tens[3] ;
 wire \u_n2a2.hundreds[0] ;
 wire \u_n2a2.hundreds[1] ;
 wire \u_n2a2.ones[0] ;
 wire \u_n2a2.ones[1] ;
 wire \u_n2a2.ones[2] ;
 wire \u_n2a2.ones[3] ;
 wire \u_n2a2.tens[0] ;
 wire \u_n2a2.tens[1] ;
 wire \u_n2a2.tens[2] ;
 wire \u_n2a2.tens[3] ;
 wire \u_n2a3.hundreds[0] ;
 wire \u_n2a3.hundreds[1] ;
 wire \u_n2a3.ones[0] ;
 wire \u_n2a3.ones[1] ;
 wire \u_n2a3.ones[2] ;
 wire \u_n2a3.ones[3] ;
 wire \u_n2a3.tens[0] ;
 wire \u_n2a3.tens[1] ;
 wire \u_n2a3.tens[2] ;
 wire \u_n2a3.tens[3] ;
 wire \u_uart.rom.addr[0] ;
 wire \u_uart.rom.addr[10] ;
 wire \u_uart.rom.addr[11] ;
 wire \u_uart.rom.addr[12] ;
 wire \u_uart.rom.addr[13] ;
 wire \u_uart.rom.addr[14] ;
 wire \u_uart.rom.addr[15] ;
 wire \u_uart.rom.addr[16] ;
 wire \u_uart.rom.addr[17] ;
 wire \u_uart.rom.addr[18] ;
 wire \u_uart.rom.addr[19] ;
 wire \u_uart.rom.addr[1] ;
 wire \u_uart.rom.addr[20] ;
 wire \u_uart.rom.addr[21] ;
 wire \u_uart.rom.addr[22] ;
 wire \u_uart.rom.addr[23] ;
 wire \u_uart.rom.addr[24] ;
 wire \u_uart.rom.addr[25] ;
 wire \u_uart.rom.addr[26] ;
 wire \u_uart.rom.addr[27] ;
 wire \u_uart.rom.addr[28] ;
 wire \u_uart.rom.addr[29] ;
 wire \u_uart.rom.addr[2] ;
 wire \u_uart.rom.addr[30] ;
 wire \u_uart.rom.addr[31] ;
 wire \u_uart.rom.addr[3] ;
 wire \u_uart.rom.addr[4] ;
 wire \u_uart.rom.addr[5] ;
 wire \u_uart.rom.addr[6] ;
 wire \u_uart.rom.addr[7] ;
 wire \u_uart.rom.addr[8] ;
 wire \u_uart.rom.addr[9] ;
 wire \u_uart.state[0] ;
 wire \u_uart.state[1] ;
 wire \u_uart.state[2] ;
 wire \u_uart.state[3] ;
 wire \u_uart.uart_tx_inst.bit_index[0] ;
 wire \u_uart.uart_tx_inst.bit_index[1] ;
 wire \u_uart.uart_tx_inst.bit_index[2] ;
 wire \u_uart.uart_tx_inst.clk_count[0] ;
 wire \u_uart.uart_tx_inst.clk_count[10] ;
 wire \u_uart.uart_tx_inst.clk_count[11] ;
 wire \u_uart.uart_tx_inst.clk_count[12] ;
 wire \u_uart.uart_tx_inst.clk_count[13] ;
 wire \u_uart.uart_tx_inst.clk_count[14] ;
 wire \u_uart.uart_tx_inst.clk_count[15] ;
 wire \u_uart.uart_tx_inst.clk_count[16] ;
 wire \u_uart.uart_tx_inst.clk_count[17] ;
 wire \u_uart.uart_tx_inst.clk_count[18] ;
 wire \u_uart.uart_tx_inst.clk_count[19] ;
 wire \u_uart.uart_tx_inst.clk_count[1] ;
 wire \u_uart.uart_tx_inst.clk_count[20] ;
 wire \u_uart.uart_tx_inst.clk_count[21] ;
 wire \u_uart.uart_tx_inst.clk_count[22] ;
 wire \u_uart.uart_tx_inst.clk_count[23] ;
 wire \u_uart.uart_tx_inst.clk_count[24] ;
 wire \u_uart.uart_tx_inst.clk_count[25] ;
 wire \u_uart.uart_tx_inst.clk_count[26] ;
 wire \u_uart.uart_tx_inst.clk_count[27] ;
 wire \u_uart.uart_tx_inst.clk_count[28] ;
 wire \u_uart.uart_tx_inst.clk_count[29] ;
 wire \u_uart.uart_tx_inst.clk_count[2] ;
 wire \u_uart.uart_tx_inst.clk_count[30] ;
 wire \u_uart.uart_tx_inst.clk_count[31] ;
 wire \u_uart.uart_tx_inst.clk_count[3] ;
 wire \u_uart.uart_tx_inst.clk_count[4] ;
 wire \u_uart.uart_tx_inst.clk_count[5] ;
 wire \u_uart.uart_tx_inst.clk_count[6] ;
 wire \u_uart.uart_tx_inst.clk_count[7] ;
 wire \u_uart.uart_tx_inst.clk_count[8] ;
 wire \u_uart.uart_tx_inst.clk_count[9] ;
 wire \u_uart.uart_tx_inst.state[0] ;
 wire \u_uart.uart_tx_inst.state[1] ;
 wire \u_uart.uart_tx_inst.state[2] ;
 wire \u_uart.uart_tx_inst.state[3] ;
 wire \u_uart.uart_tx_inst.state[4] ;
 wire \u_uart.uart_tx_inst.tx_data[0] ;
 wire \u_uart.uart_tx_inst.tx_data[1] ;
 wire \u_uart.uart_tx_inst.tx_data[2] ;
 wire \u_uart.uart_tx_inst.tx_data[3] ;
 wire \u_uart.uart_tx_inst.tx_data[4] ;
 wire \u_uart.uart_tx_inst.tx_data[5] ;
 wire \u_uart.uart_tx_inst.tx_data[6] ;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire [0:0] \u_uart.uart_tx_inst.i_Tx_Start ;

 sg13g2_inv_1 _1600_ (.Y(_0926_),
    .A(net762));
 sg13g2_inv_1 _1601_ (.Y(_0927_),
    .A(net744));
 sg13g2_inv_1 _1602_ (.Y(_0928_),
    .A(net761));
 sg13g2_inv_1 _1603_ (.Y(_0929_),
    .A(net774));
 sg13g2_inv_1 _1604_ (.Y(_0930_),
    .A(net687));
 sg13g2_inv_1 _1605_ (.Y(_0931_),
    .A(\u_uart.rom.addr[15] ));
 sg13g2_inv_1 _1606_ (.Y(_0932_),
    .A(\u_uart.rom.addr[14] ));
 sg13g2_inv_1 _1607_ (.Y(_0933_),
    .A(net611));
 sg13g2_inv_1 _1608_ (.Y(_0934_),
    .A(net637));
 sg13g2_inv_1 _1609_ (.Y(_0935_),
    .A(\u_uart.rom.addr[8] ));
 sg13g2_inv_2 _1610_ (.Y(_0936_),
    .A(net815));
 sg13g2_inv_2 _1611_ (.Y(_0937_),
    .A(net864));
 sg13g2_inv_1 _1612_ (.Y(_0938_),
    .A(net895));
 sg13g2_inv_1 _1613_ (.Y(_0939_),
    .A(\u_uart.uart_tx_inst.i_Tx_Start [0]));
 sg13g2_inv_1 _1614_ (.Y(_0940_),
    .A(o_Tx_Serial));
 sg13g2_inv_1 _1615_ (.Y(_0941_),
    .A(net564));
 sg13g2_inv_1 _1616_ (.Y(_0942_),
    .A(net562));
 sg13g2_inv_1 _1617_ (.Y(_0943_),
    .A(net152));
 sg13g2_inv_1 _1618_ (.Y(_0944_),
    .A(\u_cnt3.count[2] ));
 sg13g2_inv_1 _1619_ (.Y(_0945_),
    .A(net587));
 sg13g2_inv_2 _1620_ (.Y(_0946_),
    .A(net154));
 sg13g2_inv_2 _1621_ (.Y(_0947_),
    .A(\u_cnt2.count[3] ));
 sg13g2_inv_4 _1622_ (.A(net852),
    .Y(_0948_));
 sg13g2_inv_1 _1623_ (.Y(_0949_),
    .A(net571));
 sg13g2_inv_4 _1624_ (.A(\u_cnt1.count[4] ),
    .Y(_0950_));
 sg13g2_inv_2 _1625_ (.Y(_0951_),
    .A(net857));
 sg13g2_inv_1 _1626_ (.Y(_0952_),
    .A(net156));
 sg13g2_inv_2 _1627_ (.Y(_0953_),
    .A(net856));
 sg13g2_inv_1 _1628_ (.Y(_0954_),
    .A(net646));
 sg13g2_inv_1 _1629_ (.Y(_0955_),
    .A(net588));
 sg13g2_inv_2 _1630_ (.Y(_0956_),
    .A(net583));
 sg13g2_inv_2 _1631_ (.Y(_0957_),
    .A(net573));
 sg13g2_inv_1 _1632_ (.Y(_0958_),
    .A(net765));
 sg13g2_inv_2 _1633_ (.Y(_0959_),
    .A(net589));
 sg13g2_inv_1 _1634_ (.Y(_0960_),
    .A(net173));
 sg13g2_inv_1 _1635_ (.Y(_0961_),
    .A(net723));
 sg13g2_nor2b_1 _1636_ (.A(net802),
    .B_N(\u_uart.state[0] ),
    .Y(_0962_));
 sg13g2_or3_1 _1637_ (.A(net166),
    .B(net548),
    .C(net803),
    .X(_0002_));
 sg13g2_nand3_1 _1638_ (.B(\u_uart.uart_tx_inst.clk_count[3] ),
    .C(\u_uart.uart_tx_inst.clk_count[2] ),
    .A(net562),
    .Y(_0963_));
 sg13g2_inv_1 _1639_ (.Y(_0964_),
    .A(_0963_));
 sg13g2_nand2_1 _1640_ (.Y(_0965_),
    .A(net780),
    .B(_0964_));
 sg13g2_nor4_1 _1641_ (.A(\u_uart.uart_tx_inst.clk_count[9] ),
    .B(\u_uart.uart_tx_inst.clk_count[8] ),
    .C(\u_uart.uart_tx_inst.clk_count[7] ),
    .D(\u_uart.uart_tx_inst.clk_count[6] ),
    .Y(_0966_));
 sg13g2_a21oi_1 _1642_ (.A1(_0965_),
    .A2(_0966_),
    .Y(_0967_),
    .B1(_0941_));
 sg13g2_nor2_1 _1643_ (.A(net490),
    .B(net493),
    .Y(_0968_));
 sg13g2_nor4_1 _1644_ (.A(net506),
    .B(net492),
    .C(net481),
    .D(net475),
    .Y(_0969_));
 sg13g2_nor3_1 _1645_ (.A(net512),
    .B(net478),
    .C(net486),
    .Y(_0970_));
 sg13g2_nor4_1 _1646_ (.A(net497),
    .B(net487),
    .C(net502),
    .D(net474),
    .Y(_0971_));
 sg13g2_nor4_1 _1647_ (.A(net500),
    .B(net484),
    .C(net482),
    .D(net494),
    .Y(_0972_));
 sg13g2_nor4_1 _1648_ (.A(net488),
    .B(net479),
    .C(net498),
    .D(net476),
    .Y(_0973_));
 sg13g2_nand2_1 _1649_ (.Y(_0974_),
    .A(_0972_),
    .B(_0973_));
 sg13g2_nand4_1 _1650_ (.B(_0969_),
    .C(_0970_),
    .A(_0968_),
    .Y(_0975_),
    .D(_0971_));
 sg13g2_nor3_2 _1651_ (.A(_0967_),
    .B(_0974_),
    .C(_0975_),
    .Y(_0976_));
 sg13g2_nand2_1 _1652_ (.Y(_0977_),
    .A(net561),
    .B(_0976_));
 sg13g2_nand3_1 _1653_ (.B(net862),
    .C(\u_uart.uart_tx_inst.bit_index[0] ),
    .A(net536),
    .Y(_0978_));
 sg13g2_nor2_1 _1654_ (.A(_0976_),
    .B(net863),
    .Y(_0979_));
 sg13g2_nand2_1 _1655_ (.Y(_0980_),
    .A(net723),
    .B(_0979_));
 sg13g2_a21oi_1 _1656_ (.A1(_0977_),
    .A2(net724),
    .Y(_0008_),
    .B1(net163));
 sg13g2_nor2_1 _1657_ (.A(net163),
    .B(_0976_),
    .Y(_0981_));
 sg13g2_nor3_1 _1658_ (.A(net163),
    .B(_0961_),
    .C(_0979_),
    .Y(_0982_));
 sg13g2_a21o_1 _1659_ (.A2(_0981_),
    .A1(net850),
    .B1(_0982_),
    .X(_0006_));
 sg13g2_and2_1 _1660_ (.A(net851),
    .B(net825),
    .X(_0983_));
 sg13g2_nand2_2 _1661_ (.Y(_0984_),
    .A(\u_uart.uart_tx_inst.i_Tx_Start [0]),
    .B(\u_uart.uart_tx_inst.state[0] ));
 sg13g2_a21oi_1 _1662_ (.A1(net850),
    .A2(_0976_),
    .Y(_0985_),
    .B1(net146));
 sg13g2_nor2_1 _1663_ (.A(net163),
    .B(_0985_),
    .Y(_0007_));
 sg13g2_nand2b_1 _1664_ (.Y(_0986_),
    .B(\u_uart.state[1] ),
    .A_N(net606));
 sg13g2_nand2b_1 _1665_ (.Y(_0987_),
    .B(net714),
    .A_N(o_Tx_Active));
 sg13g2_a21oi_1 _1666_ (.A1(_0986_),
    .A2(net715),
    .Y(_0003_),
    .B1(net166));
 sg13g2_a21oi_1 _1667_ (.A1(_0939_),
    .A2(\u_uart.uart_tx_inst.state[0] ),
    .Y(_0988_),
    .B1(net164));
 sg13g2_nand2b_1 _1668_ (.Y(_0005_),
    .B(_0988_),
    .A_N(net541));
 sg13g2_nand2_2 _1669_ (.Y(_0989_),
    .A(net886),
    .B(net876));
 sg13g2_nor3_1 _1670_ (.A(net848),
    .B(net154),
    .C(net880),
    .Y(_0990_));
 sg13g2_or2_1 _1671_ (.X(_0991_),
    .B(_0990_),
    .A(_0989_));
 sg13g2_inv_1 _1672_ (.Y(_0287_),
    .A(_0991_));
 sg13g2_nor3_2 _1673_ (.A(\u_cnt2.count[3] ),
    .B(_0989_),
    .C(_0990_),
    .Y(_0992_));
 sg13g2_and2_1 _1674_ (.A(\u_cnt2.count[3] ),
    .B(_0989_),
    .X(_0993_));
 sg13g2_nor2_1 _1675_ (.A(_0992_),
    .B(_0993_),
    .Y(_0994_));
 sg13g2_nor4_1 _1676_ (.A(net154),
    .B(net852),
    .C(_0992_),
    .D(_0993_),
    .Y(_0995_));
 sg13g2_nand3_1 _1677_ (.B(_0948_),
    .C(_0994_),
    .A(_0946_),
    .Y(_0996_));
 sg13g2_nand2_1 _1678_ (.Y(_0997_),
    .A(net876),
    .B(_0991_));
 sg13g2_nand2_1 _1679_ (.Y(_0998_),
    .A(_0946_),
    .B(_0992_));
 sg13g2_nand2_1 _1680_ (.Y(_0999_),
    .A(net848),
    .B(_0998_));
 sg13g2_nand3_1 _1681_ (.B(net848),
    .C(_0989_),
    .A(net876),
    .Y(_1000_));
 sg13g2_nor2_1 _1682_ (.A(_0995_),
    .B(_1000_),
    .Y(_1001_));
 sg13g2_nand2_1 _1683_ (.Y(_1002_),
    .A(net886),
    .B(_0991_));
 sg13g2_o21ai_1 _1684_ (.B1(_1002_),
    .Y(_0286_),
    .A1(_0995_),
    .A2(_1000_));
 sg13g2_nand2b_1 _1685_ (.Y(_1003_),
    .B(\u_cnt2.count[7] ),
    .A_N(\u_cnt2.count[5] ));
 sg13g2_nor2_1 _1686_ (.A(\u_cnt2.count[6] ),
    .B(_1003_),
    .Y(_1004_));
 sg13g2_and2_1 _1687_ (.A(\u_cnt2.count[6] ),
    .B(_1003_),
    .X(_1005_));
 sg13g2_a21oi_1 _1688_ (.A1(\u_cnt2.count[7] ),
    .A2(\u_cnt2.count[6] ),
    .Y(_1006_),
    .B1(\u_cnt2.count[5] ));
 sg13g2_and2_1 _1689_ (.A(\u_cnt2.count[7] ),
    .B(\u_cnt2.count[5] ),
    .X(_1007_));
 sg13g2_nor2_1 _1690_ (.A(_1006_),
    .B(_1007_),
    .Y(_1008_));
 sg13g2_nor2_1 _1691_ (.A(net154),
    .B(_1008_),
    .Y(_1009_));
 sg13g2_o21ai_1 _1692_ (.B1(_0946_),
    .Y(_1010_),
    .A1(_1006_),
    .A2(_1007_));
 sg13g2_a21oi_1 _1693_ (.A1(_1005_),
    .A2(_1010_),
    .Y(_1011_),
    .B1(_1004_));
 sg13g2_xnor2_1 _1694_ (.Y(_1012_),
    .A(_0946_),
    .B(_1011_));
 sg13g2_o21ai_1 _1695_ (.B1(_1008_),
    .Y(_1013_),
    .A1(net154),
    .A2(_1011_));
 sg13g2_nand2_1 _1696_ (.Y(_1014_),
    .A(_0946_),
    .B(_1004_));
 sg13g2_nand2_1 _1697_ (.Y(_1015_),
    .A(_1013_),
    .B(_1014_));
 sg13g2_a22oi_1 _1698_ (.Y(_1016_),
    .B1(_1013_),
    .B2(_1014_),
    .A2(_1012_),
    .A1(_0947_));
 sg13g2_a22oi_1 _1699_ (.Y(_1017_),
    .B1(_1005_),
    .B2(_1009_),
    .A2(_1004_),
    .A1(net154));
 sg13g2_inv_1 _1700_ (.Y(_1018_),
    .A(_1017_));
 sg13g2_a21oi_1 _1701_ (.A1(_0947_),
    .A2(_1012_),
    .Y(_1019_),
    .B1(_1017_));
 sg13g2_nor2_1 _1702_ (.A(_1015_),
    .B(_1019_),
    .Y(_1020_));
 sg13g2_nor2_1 _1703_ (.A(_1016_),
    .B(_1020_),
    .Y(_1021_));
 sg13g2_o21ai_1 _1704_ (.B1(_0947_),
    .Y(_1022_),
    .A1(_1016_),
    .A2(_1018_));
 sg13g2_xor2_1 _1705_ (.B(_1022_),
    .A(_1012_),
    .X(_1023_));
 sg13g2_nand3b_1 _1706_ (.B(_1017_),
    .C(\u_cnt2.count[3] ),
    .Y(_1024_),
    .A_N(_1016_));
 sg13g2_and2_1 _1707_ (.A(_1022_),
    .B(_1024_),
    .X(_1025_));
 sg13g2_nand3_1 _1708_ (.B(_1022_),
    .C(_1024_),
    .A(_0948_),
    .Y(_1026_));
 sg13g2_a21oi_1 _1709_ (.A1(_1023_),
    .A2(_1026_),
    .Y(_1027_),
    .B1(_1021_));
 sg13g2_nor2_1 _1710_ (.A(net852),
    .B(_1027_),
    .Y(_1028_));
 sg13g2_xnor2_1 _1711_ (.Y(_1029_),
    .A(_0948_),
    .B(_1027_));
 sg13g2_and2_1 _1712_ (.A(_0949_),
    .B(_1029_),
    .X(_1030_));
 sg13g2_xnor2_1 _1713_ (.Y(_1031_),
    .A(_1025_),
    .B(_1028_));
 sg13g2_nand2b_1 _1714_ (.Y(_1032_),
    .B(_1031_),
    .A_N(_1030_));
 sg13g2_and3_2 _1715_ (.X(_1033_),
    .A(_0947_),
    .B(_0948_),
    .C(_0286_));
 sg13g2_a21oi_1 _1716_ (.A1(_0948_),
    .A2(_0286_),
    .Y(_1034_),
    .B1(_0994_));
 sg13g2_nor2_2 _1717_ (.A(_1033_),
    .B(_1034_),
    .Y(_1035_));
 sg13g2_nand2_1 _1718_ (.Y(_1036_),
    .A(_0996_),
    .B(_0286_));
 sg13g2_nand3b_1 _1719_ (.B(_0286_),
    .C(_0996_),
    .Y(_1037_),
    .A_N(_0999_));
 sg13g2_xor2_1 _1720_ (.B(_1036_),
    .A(_0999_),
    .X(_1038_));
 sg13g2_xnor2_1 _1721_ (.Y(_1039_),
    .A(\u_cnt2.count[4] ),
    .B(_0992_));
 sg13g2_xnor2_1 _1722_ (.Y(_1040_),
    .A(_1033_),
    .B(_1039_));
 sg13g2_a21oi_1 _1723_ (.A1(_0997_),
    .A2(_1037_),
    .Y(_1041_),
    .B1(_1001_));
 sg13g2_a21o_1 _1724_ (.A2(_1037_),
    .A1(_0997_),
    .B1(_1001_),
    .X(_1042_));
 sg13g2_o21ai_1 _1725_ (.B1(_1041_),
    .Y(_1043_),
    .A1(_1038_),
    .A2(_1040_));
 sg13g2_inv_1 _1726_ (.Y(_0291_),
    .A(_1043_));
 sg13g2_nand3b_1 _1727_ (.B(_1041_),
    .C(_1038_),
    .Y(_1044_),
    .A_N(_1040_));
 sg13g2_and2_1 _1728_ (.A(_1038_),
    .B(_1044_),
    .X(_1045_));
 sg13g2_nand2_1 _1729_ (.Y(_1046_),
    .A(_1040_),
    .B(_1042_));
 sg13g2_nand2_1 _1730_ (.Y(_1047_),
    .A(_1044_),
    .B(_1046_));
 sg13g2_nand3_1 _1731_ (.B(_1044_),
    .C(_1046_),
    .A(_1035_),
    .Y(_1048_));
 sg13g2_nor3_1 _1732_ (.A(_1038_),
    .B(_1040_),
    .C(_1042_),
    .Y(_1049_));
 sg13g2_a21oi_1 _1733_ (.A1(_1045_),
    .A2(_1048_),
    .Y(_1050_),
    .B1(_1049_));
 sg13g2_inv_1 _1734_ (.Y(_0290_),
    .A(_1050_));
 sg13g2_xnor2_1 _1735_ (.Y(_1051_),
    .A(_0948_),
    .B(_0286_));
 sg13g2_xnor2_1 _1736_ (.Y(_1052_),
    .A(_1035_),
    .B(_1050_));
 sg13g2_xnor2_1 _1737_ (.Y(_1053_),
    .A(_1035_),
    .B(_0290_));
 sg13g2_a21oi_1 _1738_ (.A1(_1035_),
    .A2(_1049_),
    .Y(_1054_),
    .B1(_1047_));
 sg13g2_nand4_1 _1739_ (.B(_1038_),
    .C(_1040_),
    .A(_1035_),
    .Y(_1055_),
    .D(_1042_));
 sg13g2_nor2b_1 _1740_ (.A(_1054_),
    .B_N(_1055_),
    .Y(_1056_));
 sg13g2_a21oi_1 _1741_ (.A1(_1048_),
    .A2(_1049_),
    .Y(_1057_),
    .B1(_1045_));
 sg13g2_a21oi_1 _1742_ (.A1(_1045_),
    .A2(_1048_),
    .Y(_1058_),
    .B1(_1057_));
 sg13g2_o21ai_1 _1743_ (.B1(_1058_),
    .Y(_1059_),
    .A1(_1051_),
    .A2(_1053_));
 sg13g2_nand3b_1 _1744_ (.B(_1052_),
    .C(_1056_),
    .Y(_1060_),
    .A_N(_1051_));
 sg13g2_nand2_1 _1745_ (.Y(_1061_),
    .A(_1059_),
    .B(_1060_));
 sg13g2_nand3_1 _1746_ (.B(_1059_),
    .C(_1060_),
    .A(_1032_),
    .Y(_0288_));
 sg13g2_o21ai_1 _1747_ (.B1(_1056_),
    .Y(_1062_),
    .A1(_1051_),
    .A2(_1053_));
 sg13g2_nand2b_1 _1748_ (.Y(_0289_),
    .B(_1062_),
    .A_N(_1058_));
 sg13g2_nand2b_2 _1749_ (.Y(_1063_),
    .B(\u_uart.rom.addr[0] ),
    .A_N(\u_uart.rom.addr[1] ));
 sg13g2_nand2b_2 _1750_ (.Y(_1064_),
    .B(net147),
    .A_N(net149));
 sg13g2_nor2_1 _1751_ (.A(_1063_),
    .B(_1064_),
    .Y(_1065_));
 sg13g2_nor2_1 _1752_ (.A(\u_uart.rom.addr[7] ),
    .B(\u_uart.rom.addr[6] ),
    .Y(_1066_));
 sg13g2_nand3_1 _1753_ (.B(_0937_),
    .C(_1066_),
    .A(\u_uart.rom.addr[5] ),
    .Y(_1067_));
 sg13g2_nor4_1 _1754_ (.A(\u_uart.rom.addr[27] ),
    .B(\u_uart.rom.addr[26] ),
    .C(\u_uart.rom.addr[25] ),
    .D(\u_uart.rom.addr[24] ),
    .Y(_1068_));
 sg13g2_nor4_1 _1755_ (.A(\u_uart.rom.addr[31] ),
    .B(\u_uart.rom.addr[30] ),
    .C(\u_uart.rom.addr[29] ),
    .D(\u_uart.rom.addr[28] ),
    .Y(_1069_));
 sg13g2_nand2_1 _1756_ (.Y(_1070_),
    .A(_1068_),
    .B(_1069_));
 sg13g2_nor4_1 _1757_ (.A(\u_uart.rom.addr[19] ),
    .B(\u_uart.rom.addr[18] ),
    .C(\u_uart.rom.addr[17] ),
    .D(\u_uart.rom.addr[16] ),
    .Y(_1071_));
 sg13g2_nor4_1 _1758_ (.A(\u_uart.rom.addr[23] ),
    .B(\u_uart.rom.addr[22] ),
    .C(\u_uart.rom.addr[21] ),
    .D(\u_uart.rom.addr[20] ),
    .Y(_1072_));
 sg13g2_nor4_1 _1759_ (.A(\u_uart.rom.addr[11] ),
    .B(\u_uart.rom.addr[10] ),
    .C(\u_uart.rom.addr[9] ),
    .D(\u_uart.rom.addr[8] ),
    .Y(_1073_));
 sg13g2_or4_1 _1760_ (.A(\u_uart.rom.addr[15] ),
    .B(\u_uart.rom.addr[14] ),
    .C(\u_uart.rom.addr[13] ),
    .D(\u_uart.rom.addr[12] ),
    .X(_1074_));
 sg13g2_nand3_1 _1761_ (.B(_1072_),
    .C(_1073_),
    .A(_1071_),
    .Y(_1075_));
 sg13g2_nor3_2 _1762_ (.A(_1070_),
    .B(_1074_),
    .C(_1075_),
    .Y(_1076_));
 sg13g2_nor2b_2 _1763_ (.A(_1067_),
    .B_N(_1076_),
    .Y(_1077_));
 sg13g2_inv_1 _1764_ (.Y(_1078_),
    .A(_1077_));
 sg13g2_and2_1 _1765_ (.A(_1065_),
    .B(_1077_),
    .X(_1079_));
 sg13g2_nand2_1 _1766_ (.Y(_1080_),
    .A(_1065_),
    .B(_1077_));
 sg13g2_nand3_1 _1767_ (.B(net846),
    .C(_1080_),
    .A(net606),
    .Y(_1081_));
 sg13g2_nand2_1 _1768_ (.Y(_1082_),
    .A(o_Tx_Active),
    .B(\u_uart.state[2] ));
 sg13g2_a22oi_1 _1769_ (.Y(_1083_),
    .B1(net714),
    .B2(net728),
    .A2(\u_uart.state[0] ),
    .A1(net802));
 sg13g2_a21oi_1 _1770_ (.A1(_1081_),
    .A2(_1083_),
    .Y(_0004_),
    .B1(net166));
 sg13g2_nand2_2 _1771_ (.Y(_1084_),
    .A(net888),
    .B(net151));
 sg13g2_nor3_1 _1772_ (.A(net870),
    .B(net152),
    .C(net153),
    .Y(_1085_));
 sg13g2_or2_1 _1773_ (.X(_1086_),
    .B(_1085_),
    .A(_1084_));
 sg13g2_inv_1 _1774_ (.Y(_0296_),
    .A(_1086_));
 sg13g2_nor3_2 _1775_ (.A(net153),
    .B(_1084_),
    .C(_1085_),
    .Y(_1087_));
 sg13g2_and2_1 _1776_ (.A(net153),
    .B(_1084_),
    .X(_1088_));
 sg13g2_nor2_1 _1777_ (.A(_1087_),
    .B(_1088_),
    .Y(_1089_));
 sg13g2_nor4_1 _1778_ (.A(net152),
    .B(net894),
    .C(_1087_),
    .D(_1088_),
    .Y(_1090_));
 sg13g2_nand2_1 _1779_ (.Y(_1091_),
    .A(_0943_),
    .B(_1087_));
 sg13g2_nand2_1 _1780_ (.Y(_1092_),
    .A(net902),
    .B(_1091_));
 sg13g2_nand3_1 _1781_ (.B(net870),
    .C(_1084_),
    .A(net151),
    .Y(_1093_));
 sg13g2_nor2_1 _1782_ (.A(_1090_),
    .B(_1092_),
    .Y(_1094_));
 sg13g2_nor2_1 _1783_ (.A(_1090_),
    .B(_1093_),
    .Y(_1095_));
 sg13g2_nand2_1 _1784_ (.Y(_1096_),
    .A(net888),
    .B(_1086_));
 sg13g2_o21ai_1 _1785_ (.B1(_1096_),
    .Y(_0295_),
    .A1(_1090_),
    .A2(_1093_));
 sg13g2_nand2b_1 _1786_ (.Y(_1097_),
    .B(\u_cnt3.count[7] ),
    .A_N(\u_cnt3.count[5] ));
 sg13g2_nor2_1 _1787_ (.A(net151),
    .B(_1097_),
    .Y(_1098_));
 sg13g2_and2_1 _1788_ (.A(\u_cnt3.count[6] ),
    .B(_1097_),
    .X(_1099_));
 sg13g2_nand2_1 _1789_ (.Y(_1100_),
    .A(net151),
    .B(_1097_));
 sg13g2_a21oi_1 _1790_ (.A1(\u_cnt3.count[7] ),
    .A2(net151),
    .Y(_1101_),
    .B1(\u_cnt3.count[5] ));
 sg13g2_and2_1 _1791_ (.A(\u_cnt3.count[7] ),
    .B(\u_cnt3.count[5] ),
    .X(_1102_));
 sg13g2_nor2_1 _1792_ (.A(_1101_),
    .B(_1102_),
    .Y(_1103_));
 sg13g2_o21ai_1 _1793_ (.B1(_0943_),
    .Y(_1104_),
    .A1(_1101_),
    .A2(_1102_));
 sg13g2_a21oi_1 _1794_ (.A1(_1099_),
    .A2(_1104_),
    .Y(_1105_),
    .B1(_1098_));
 sg13g2_xnor2_1 _1795_ (.Y(_1106_),
    .A(net152),
    .B(_1105_));
 sg13g2_or2_1 _1796_ (.X(_1107_),
    .B(_1106_),
    .A(net153));
 sg13g2_nand2_1 _1797_ (.Y(_1108_),
    .A(_0943_),
    .B(_1098_));
 sg13g2_o21ai_1 _1798_ (.B1(_1103_),
    .Y(_1109_),
    .A1(net152),
    .A2(_1105_));
 sg13g2_nand2_1 _1799_ (.Y(_1110_),
    .A(_1108_),
    .B(_1109_));
 sg13g2_nand2_1 _1800_ (.Y(_1111_),
    .A(net152),
    .B(_1098_));
 sg13g2_o21ai_1 _1801_ (.B1(_1111_),
    .Y(_1112_),
    .A1(_1100_),
    .A2(_1104_));
 sg13g2_a21oi_1 _1802_ (.A1(_1107_),
    .A2(_1110_),
    .Y(_1113_),
    .B1(_1112_));
 sg13g2_nor2_1 _1803_ (.A(\u_cnt3.count[3] ),
    .B(_1113_),
    .Y(_1114_));
 sg13g2_xnor2_1 _1804_ (.Y(_1115_),
    .A(net153),
    .B(_1113_));
 sg13g2_inv_1 _1805_ (.Y(_1116_),
    .A(_1115_));
 sg13g2_a21oi_1 _1806_ (.A1(_1107_),
    .A2(_1112_),
    .Y(_1117_),
    .B1(_1110_));
 sg13g2_a21oi_1 _1807_ (.A1(_1107_),
    .A2(_1110_),
    .Y(_1118_),
    .B1(_1117_));
 sg13g2_nand2b_1 _1808_ (.Y(_1119_),
    .B(_0944_),
    .A_N(_1115_));
 sg13g2_xor2_1 _1809_ (.B(_1114_),
    .A(_1106_),
    .X(_1120_));
 sg13g2_a21oi_2 _1810_ (.B1(_1118_),
    .Y(_1121_),
    .A2(_1120_),
    .A1(_1119_));
 sg13g2_nand2_1 _1811_ (.Y(_1122_),
    .A(net875),
    .B(_1121_));
 sg13g2_a21oi_1 _1812_ (.A1(_1120_),
    .A2(_1121_),
    .Y(_1123_),
    .B1(_1118_));
 sg13g2_nor2_1 _1813_ (.A(net875),
    .B(_1121_),
    .Y(_1124_));
 sg13g2_o21ai_1 _1814_ (.B1(_1123_),
    .Y(_1125_),
    .A1(_1116_),
    .A2(_1122_));
 sg13g2_xnor2_1 _1815_ (.Y(_1126_),
    .A(net875),
    .B(_1121_));
 sg13g2_nor3_1 _1816_ (.A(_0945_),
    .B(_1116_),
    .C(_1126_),
    .Y(_1127_));
 sg13g2_nor2_2 _1817_ (.A(_1125_),
    .B(_1127_),
    .Y(_1128_));
 sg13g2_inv_1 _1818_ (.Y(_0297_),
    .A(_1128_));
 sg13g2_a21oi_1 _1819_ (.A1(_1093_),
    .A2(_1096_),
    .Y(_1129_),
    .B1(_1090_));
 sg13g2_xnor2_1 _1820_ (.Y(_1130_),
    .A(_1092_),
    .B(_1129_));
 sg13g2_and2_1 _1821_ (.A(_0944_),
    .B(_0295_),
    .X(_1131_));
 sg13g2_nor2b_1 _1822_ (.A(net153),
    .B_N(_1131_),
    .Y(_1132_));
 sg13g2_xnor2_1 _1823_ (.Y(_1133_),
    .A(net152),
    .B(_1087_));
 sg13g2_xnor2_1 _1824_ (.Y(_1134_),
    .A(_1132_),
    .B(_1133_));
 sg13g2_a22oi_1 _1825_ (.Y(_1135_),
    .B1(_1094_),
    .B2(_0295_),
    .A2(_1086_),
    .A1(net151));
 sg13g2_or2_1 _1826_ (.X(_1136_),
    .B(_1135_),
    .A(_1095_));
 sg13g2_nor2_1 _1827_ (.A(_1134_),
    .B(_1136_),
    .Y(_1137_));
 sg13g2_nor2_1 _1828_ (.A(_1089_),
    .B(_1131_),
    .Y(_1138_));
 sg13g2_nor2_1 _1829_ (.A(_1132_),
    .B(_1138_),
    .Y(_1139_));
 sg13g2_and2_1 _1830_ (.A(_1134_),
    .B(_1136_),
    .X(_1140_));
 sg13g2_nor2_1 _1831_ (.A(_1130_),
    .B(_1134_),
    .Y(_1141_));
 sg13g2_nor2_1 _1832_ (.A(_1136_),
    .B(_1141_),
    .Y(_0300_));
 sg13g2_a21oi_1 _1833_ (.A1(_1130_),
    .A2(_1137_),
    .Y(_1142_),
    .B1(_1140_));
 sg13g2_and2_1 _1834_ (.A(_1139_),
    .B(_1142_),
    .X(_1143_));
 sg13g2_nor2b_1 _1835_ (.A(_1137_),
    .B_N(_1130_),
    .Y(_1144_));
 sg13g2_nand2_1 _1836_ (.Y(_1145_),
    .A(_1143_),
    .B(_1144_));
 sg13g2_nor3_1 _1837_ (.A(_1130_),
    .B(_1134_),
    .C(_1136_),
    .Y(_1146_));
 sg13g2_nor2b_1 _1838_ (.A(_1143_),
    .B_N(_1144_),
    .Y(_1147_));
 sg13g2_or2_1 _1839_ (.X(_0299_),
    .B(_1147_),
    .A(_1146_));
 sg13g2_nor2_1 _1840_ (.A(_0944_),
    .B(_0295_),
    .Y(_1148_));
 sg13g2_nor3_1 _1841_ (.A(_1131_),
    .B(_1146_),
    .C(_1148_),
    .Y(_1149_));
 sg13g2_and2_1 _1842_ (.A(_0299_),
    .B(_1149_),
    .X(_1150_));
 sg13g2_o21ai_1 _1843_ (.B1(_1139_),
    .Y(_1151_),
    .A1(_1147_),
    .A2(_1149_));
 sg13g2_o21ai_1 _1844_ (.B1(_1151_),
    .Y(_1152_),
    .A1(_1137_),
    .A2(_1140_));
 sg13g2_o21ai_1 _1845_ (.B1(_1145_),
    .Y(_0298_),
    .A1(_1150_),
    .A2(_1152_));
 sg13g2_nand2_1 _1846_ (.Y(_1153_),
    .A(net878),
    .B(net853));
 sg13g2_nor3_1 _1847_ (.A(net860),
    .B(net887),
    .C(net155),
    .Y(_1154_));
 sg13g2_or2_1 _1848_ (.X(_1155_),
    .B(_1154_),
    .A(_1153_));
 sg13g2_inv_1 _1849_ (.Y(_0278_),
    .A(_1155_));
 sg13g2_nor2_2 _1850_ (.A(net155),
    .B(_1155_),
    .Y(_1156_));
 sg13g2_and2_1 _1851_ (.A(net155),
    .B(_1153_),
    .X(_1157_));
 sg13g2_nor2_1 _1852_ (.A(_1156_),
    .B(_1157_),
    .Y(_1158_));
 sg13g2_nor4_1 _1853_ (.A(\u_cnt1.count[4] ),
    .B(net882),
    .C(_1156_),
    .D(_1157_),
    .Y(_1159_));
 sg13g2_nand3_1 _1854_ (.B(_0951_),
    .C(_1158_),
    .A(_0950_),
    .Y(_1160_));
 sg13g2_nand2_1 _1855_ (.Y(_1161_),
    .A(net853),
    .B(_1155_));
 sg13g2_nand2_1 _1856_ (.Y(_1162_),
    .A(_0950_),
    .B(_1156_));
 sg13g2_nand2_1 _1857_ (.Y(_1163_),
    .A(net901),
    .B(_1162_));
 sg13g2_nand3_1 _1858_ (.B(net860),
    .C(_1153_),
    .A(net853),
    .Y(_1164_));
 sg13g2_nor2_1 _1859_ (.A(_1159_),
    .B(_1164_),
    .Y(_1165_));
 sg13g2_nand2_1 _1860_ (.Y(_1166_),
    .A(net878),
    .B(_1155_));
 sg13g2_o21ai_1 _1861_ (.B1(_1166_),
    .Y(_0277_),
    .A1(_1159_),
    .A2(_1164_));
 sg13g2_nand2b_1 _1862_ (.Y(_1167_),
    .B(\u_cnt1.count[7] ),
    .A_N(\u_cnt1.count[5] ));
 sg13g2_and2_1 _1863_ (.A(\u_cnt1.count[6] ),
    .B(_1167_),
    .X(_1168_));
 sg13g2_a21oi_1 _1864_ (.A1(\u_cnt1.count[7] ),
    .A2(\u_cnt1.count[6] ),
    .Y(_1169_),
    .B1(\u_cnt1.count[5] ));
 sg13g2_and2_1 _1865_ (.A(\u_cnt1.count[7] ),
    .B(\u_cnt1.count[5] ),
    .X(_1170_));
 sg13g2_nor2_1 _1866_ (.A(_1169_),
    .B(_1170_),
    .Y(_1171_));
 sg13g2_nor2_1 _1867_ (.A(\u_cnt1.count[4] ),
    .B(_1171_),
    .Y(_1172_));
 sg13g2_o21ai_1 _1868_ (.B1(_0950_),
    .Y(_1173_),
    .A1(_1169_),
    .A2(_1170_));
 sg13g2_nor2_1 _1869_ (.A(\u_cnt1.count[6] ),
    .B(_1167_),
    .Y(_1174_));
 sg13g2_a22oi_1 _1870_ (.Y(_1175_),
    .B1(_1174_),
    .B2(\u_cnt1.count[4] ),
    .A2(_1172_),
    .A1(_1168_));
 sg13g2_a21oi_1 _1871_ (.A1(_1168_),
    .A2(_1173_),
    .Y(_1176_),
    .B1(_1174_));
 sg13g2_or2_1 _1872_ (.X(_1177_),
    .B(_1176_),
    .A(\u_cnt1.count[4] ));
 sg13g2_xnor2_1 _1873_ (.Y(_1178_),
    .A(_0950_),
    .B(_1176_));
 sg13g2_nor2b_2 _1874_ (.A(net155),
    .B_N(_1178_),
    .Y(_1179_));
 sg13g2_a22oi_1 _1875_ (.Y(_1180_),
    .B1(_1177_),
    .B2(_1171_),
    .A2(_1174_),
    .A1(_0950_));
 sg13g2_o21ai_1 _1876_ (.B1(_1175_),
    .Y(_1181_),
    .A1(_1179_),
    .A2(_1180_));
 sg13g2_nand3_1 _1877_ (.B(_1175_),
    .C(_1180_),
    .A(net155),
    .Y(_1182_));
 sg13g2_nor2b_1 _1878_ (.A(net155),
    .B_N(_1181_),
    .Y(_1183_));
 sg13g2_xor2_1 _1879_ (.B(_1181_),
    .A(net799),
    .X(_1184_));
 sg13g2_nand2b_1 _1880_ (.Y(_1185_),
    .B(_1179_),
    .A_N(_1180_));
 sg13g2_o21ai_1 _1881_ (.B1(_1185_),
    .Y(_1186_),
    .A1(_1175_),
    .A2(_1179_));
 sg13g2_nand2b_1 _1882_ (.Y(_1187_),
    .B(_0951_),
    .A_N(_1184_));
 sg13g2_nand2b_1 _1883_ (.Y(_1188_),
    .B(_1179_),
    .A_N(_1175_));
 sg13g2_o21ai_1 _1884_ (.B1(_1188_),
    .Y(_1189_),
    .A1(_1178_),
    .A2(_1183_));
 sg13g2_a21o_1 _1885_ (.A2(_1189_),
    .A1(_1187_),
    .B1(_1186_),
    .X(_1190_));
 sg13g2_inv_1 _1886_ (.Y(_1191_),
    .A(_1190_));
 sg13g2_o21ai_1 _1887_ (.B1(_1184_),
    .Y(_1192_),
    .A1(net857),
    .A2(_1191_));
 sg13g2_xnor2_1 _1888_ (.Y(_1193_),
    .A(_0951_),
    .B(_1190_));
 sg13g2_nand2_1 _1889_ (.Y(_1194_),
    .A(net595),
    .B(_1184_));
 sg13g2_nor2_1 _1890_ (.A(_1193_),
    .B(_1194_),
    .Y(_1195_));
 sg13g2_o21ai_1 _1891_ (.B1(net857),
    .Y(_1196_),
    .A1(_1178_),
    .A2(_1183_));
 sg13g2_a22oi_1 _1892_ (.Y(_1197_),
    .B1(_1187_),
    .B2(_1196_),
    .A2(_1182_),
    .A1(_1178_));
 sg13g2_nor3_1 _1893_ (.A(_1186_),
    .B(_1195_),
    .C(_1197_),
    .Y(_1198_));
 sg13g2_inv_1 _1894_ (.Y(_0279_),
    .A(_1198_));
 sg13g2_nand2_1 _1895_ (.Y(_1199_),
    .A(_1160_),
    .B(_0277_));
 sg13g2_nand3b_1 _1896_ (.B(_0277_),
    .C(_1160_),
    .Y(_1200_),
    .A_N(_1163_));
 sg13g2_a21oi_1 _1897_ (.A1(_1161_),
    .A2(_1200_),
    .Y(_1201_),
    .B1(_1165_));
 sg13g2_xor2_1 _1898_ (.B(_1199_),
    .A(_1163_),
    .X(_1202_));
 sg13g2_and2_1 _1899_ (.A(_0951_),
    .B(_0277_),
    .X(_1203_));
 sg13g2_nand3b_1 _1900_ (.B(_0951_),
    .C(_0277_),
    .Y(_1204_),
    .A_N(net155));
 sg13g2_xnor2_1 _1901_ (.Y(_1205_),
    .A(_0950_),
    .B(_1156_));
 sg13g2_xnor2_1 _1902_ (.Y(_1206_),
    .A(_1204_),
    .B(_1205_));
 sg13g2_o21ai_1 _1903_ (.B1(_1201_),
    .Y(_1207_),
    .A1(_1202_),
    .A2(_1206_));
 sg13g2_inv_1 _1904_ (.Y(_0282_),
    .A(_1207_));
 sg13g2_and2_1 _1905_ (.A(_1201_),
    .B(_1207_),
    .X(_1208_));
 sg13g2_o21ai_1 _1906_ (.B1(_1204_),
    .Y(_1209_),
    .A1(_1158_),
    .A2(_1203_));
 sg13g2_inv_1 _1907_ (.Y(_1210_),
    .A(_1209_));
 sg13g2_a21oi_1 _1908_ (.A1(_1202_),
    .A2(_1210_),
    .Y(_1211_),
    .B1(_1208_));
 sg13g2_xor2_1 _1909_ (.B(_1207_),
    .A(_1206_),
    .X(_1212_));
 sg13g2_nor2_1 _1910_ (.A(_1209_),
    .B(_1212_),
    .Y(_1213_));
 sg13g2_o21ai_1 _1911_ (.B1(_1202_),
    .Y(_1214_),
    .A1(_1206_),
    .A2(_1207_));
 sg13g2_a21oi_1 _1912_ (.A1(_1210_),
    .A2(_1212_),
    .Y(_1215_),
    .B1(_1214_));
 sg13g2_or2_1 _1913_ (.X(_0281_),
    .B(_1215_),
    .A(_1208_));
 sg13g2_xnor2_1 _1914_ (.Y(_1216_),
    .A(net857),
    .B(_0277_));
 sg13g2_o21ai_1 _1915_ (.B1(_0281_),
    .Y(_1217_),
    .A1(_1210_),
    .A2(_1216_));
 sg13g2_a21oi_1 _1916_ (.A1(_1210_),
    .A2(_1216_),
    .Y(_1218_),
    .B1(_1212_));
 sg13g2_nand2_1 _1917_ (.Y(_1219_),
    .A(_1217_),
    .B(_1218_));
 sg13g2_o21ai_1 _1918_ (.B1(_1219_),
    .Y(_0280_),
    .A1(_1211_),
    .A2(_1213_));
 sg13g2_nand2_2 _1919_ (.Y(_1220_),
    .A(net885),
    .B(net873));
 sg13g2_nor3_1 _1920_ (.A(net869),
    .B(net156),
    .C(net874),
    .Y(_1221_));
 sg13g2_or2_1 _1921_ (.X(_1222_),
    .B(_1221_),
    .A(_1220_));
 sg13g2_inv_1 _1922_ (.Y(_0269_),
    .A(_1222_));
 sg13g2_nor3_2 _1923_ (.A(\u_cnt0.count[3] ),
    .B(_1220_),
    .C(_1221_),
    .Y(_1223_));
 sg13g2_and2_1 _1924_ (.A(\u_cnt0.count[3] ),
    .B(_1220_),
    .X(_1224_));
 sg13g2_nor2_1 _1925_ (.A(_1223_),
    .B(_1224_),
    .Y(_1225_));
 sg13g2_nor4_1 _1926_ (.A(net156),
    .B(\u_cnt0.count[2] ),
    .C(_1223_),
    .D(_1224_),
    .Y(_1226_));
 sg13g2_nand3_1 _1927_ (.B(_0953_),
    .C(_1225_),
    .A(_0952_),
    .Y(_1227_));
 sg13g2_nand2_1 _1928_ (.Y(_1228_),
    .A(net903),
    .B(_1222_));
 sg13g2_nand2_1 _1929_ (.Y(_1229_),
    .A(_0952_),
    .B(_1223_));
 sg13g2_nand2_1 _1930_ (.Y(_1230_),
    .A(\u_cnt0.count[5] ),
    .B(_1229_));
 sg13g2_nand3_1 _1931_ (.B(net869),
    .C(_1220_),
    .A(net873),
    .Y(_1231_));
 sg13g2_nor2_1 _1932_ (.A(_1226_),
    .B(_1231_),
    .Y(_1232_));
 sg13g2_nand2_1 _1933_ (.Y(_1233_),
    .A(net885),
    .B(_1222_));
 sg13g2_o21ai_1 _1934_ (.B1(_1233_),
    .Y(_0268_),
    .A1(_1226_),
    .A2(_1231_));
 sg13g2_nand2_1 _1935_ (.Y(_1234_),
    .A(_1227_),
    .B(_0268_));
 sg13g2_nand3b_1 _1936_ (.B(_0268_),
    .C(_1227_),
    .Y(_1235_),
    .A_N(_1230_));
 sg13g2_xor2_1 _1937_ (.B(_1234_),
    .A(_1230_),
    .X(_1236_));
 sg13g2_and3_2 _1938_ (.X(_1237_),
    .A(_0953_),
    .B(_1225_),
    .C(_0268_));
 sg13g2_xnor2_1 _1939_ (.Y(_1238_),
    .A(net156),
    .B(_1223_));
 sg13g2_xnor2_1 _1940_ (.Y(_1239_),
    .A(_1237_),
    .B(_1238_));
 sg13g2_a21oi_1 _1941_ (.A1(_1228_),
    .A2(_1235_),
    .Y(_1240_),
    .B1(_1232_));
 sg13g2_a21o_1 _1942_ (.A2(_1235_),
    .A1(_1228_),
    .B1(_1232_),
    .X(_1241_));
 sg13g2_o21ai_1 _1943_ (.B1(_1240_),
    .Y(_1242_),
    .A1(_1236_),
    .A2(_1239_));
 sg13g2_inv_1 _1944_ (.Y(_0273_),
    .A(_1242_));
 sg13g2_nand3b_1 _1945_ (.B(_1240_),
    .C(_1236_),
    .Y(_1243_),
    .A_N(_1239_));
 sg13g2_and2_1 _1946_ (.A(_1236_),
    .B(_1243_),
    .X(_1244_));
 sg13g2_nand2_1 _1947_ (.Y(_1245_),
    .A(_1236_),
    .B(_1243_));
 sg13g2_xnor2_1 _1948_ (.Y(_1246_),
    .A(_1239_),
    .B(_1242_));
 sg13g2_a21oi_1 _1949_ (.A1(_0953_),
    .A2(_0268_),
    .Y(_1247_),
    .B1(_1225_));
 sg13g2_nor2_2 _1950_ (.A(_1237_),
    .B(_1247_),
    .Y(_1248_));
 sg13g2_inv_1 _1951_ (.Y(_1249_),
    .A(_1248_));
 sg13g2_o21ai_1 _1952_ (.B1(_1244_),
    .Y(_1250_),
    .A1(_1246_),
    .A2(_1249_));
 sg13g2_nor3_1 _1953_ (.A(_1236_),
    .B(_1239_),
    .C(_1241_),
    .Y(_1251_));
 sg13g2_nand2_1 _1954_ (.Y(_1252_),
    .A(_1240_),
    .B(_1242_));
 sg13g2_nand2_1 _1955_ (.Y(_0272_),
    .A(_1250_),
    .B(_1252_));
 sg13g2_o21ai_1 _1956_ (.B1(_1245_),
    .Y(_1253_),
    .A1(_1248_),
    .A2(_1252_));
 sg13g2_and2_1 _1957_ (.A(_1250_),
    .B(_1253_),
    .X(_1254_));
 sg13g2_nand2_1 _1958_ (.Y(_1255_),
    .A(_1250_),
    .B(_1253_));
 sg13g2_xnor2_1 _1959_ (.Y(_1256_),
    .A(\u_cnt0.count[2] ),
    .B(_0268_));
 sg13g2_inv_1 _1960_ (.Y(_1257_),
    .A(_1256_));
 sg13g2_a221oi_1 _1961_ (.B2(_1246_),
    .C1(_1249_),
    .B1(_1244_),
    .A1(_1240_),
    .Y(_1258_),
    .A2(_1242_));
 sg13g2_a21oi_1 _1962_ (.A1(_1245_),
    .A2(_1252_),
    .Y(_1259_),
    .B1(_1248_));
 sg13g2_or2_1 _1963_ (.X(_1260_),
    .B(_1259_),
    .A(_1258_));
 sg13g2_o21ai_1 _1964_ (.B1(_1256_),
    .Y(_1261_),
    .A1(_1258_),
    .A2(_1259_));
 sg13g2_a21oi_1 _1965_ (.A1(_1248_),
    .A2(_1251_),
    .Y(_1262_),
    .B1(_1246_));
 sg13g2_nand4_1 _1966_ (.B(_1239_),
    .C(_1241_),
    .A(_1236_),
    .Y(_1263_),
    .D(_1248_));
 sg13g2_nand2b_1 _1967_ (.Y(_1264_),
    .B(_1263_),
    .A_N(_1262_));
 sg13g2_nor2b_1 _1968_ (.A(_1262_),
    .B_N(_1263_),
    .Y(_1265_));
 sg13g2_nand2_1 _1969_ (.Y(_1266_),
    .A(_1261_),
    .B(_1265_));
 sg13g2_o21ai_1 _1970_ (.B1(_1264_),
    .Y(_1267_),
    .A1(_1256_),
    .A2(_1260_));
 sg13g2_a21oi_1 _1971_ (.A1(_1266_),
    .A2(_1267_),
    .Y(_1268_),
    .B1(_1254_));
 sg13g2_a21o_1 _1972_ (.A2(_1267_),
    .A1(_1266_),
    .B1(_1254_),
    .X(_1269_));
 sg13g2_nand2_1 _1973_ (.Y(_0271_),
    .A(_1255_),
    .B(_1266_));
 sg13g2_a21oi_1 _1974_ (.A1(_1255_),
    .A2(_1264_),
    .Y(_1270_),
    .B1(_1256_));
 sg13g2_a221oi_1 _1975_ (.B2(_1265_),
    .C1(_1257_),
    .B1(_1261_),
    .A1(_1250_),
    .Y(_1271_),
    .A2(_1253_));
 sg13g2_or2_1 _1976_ (.X(_1272_),
    .B(_1271_),
    .A(_1270_));
 sg13g2_nand2b_1 _1977_ (.Y(_1273_),
    .B(\u_cnt0.count[7] ),
    .A_N(\u_cnt0.count[5] ));
 sg13g2_and2_1 _1978_ (.A(\u_cnt0.count[6] ),
    .B(_1273_),
    .X(_1274_));
 sg13g2_a21oi_1 _1979_ (.A1(\u_cnt0.count[7] ),
    .A2(\u_cnt0.count[6] ),
    .Y(_1275_),
    .B1(\u_cnt0.count[5] ));
 sg13g2_a21oi_1 _1980_ (.A1(\u_cnt0.count[7] ),
    .A2(\u_cnt0.count[5] ),
    .Y(_0304_),
    .B1(_1275_));
 sg13g2_nor2_1 _1981_ (.A(net156),
    .B(_0304_),
    .Y(_0305_));
 sg13g2_nor2_1 _1982_ (.A(\u_cnt0.count[6] ),
    .B(_1273_),
    .Y(_0306_));
 sg13g2_a22oi_1 _1983_ (.Y(_0307_),
    .B1(_0306_),
    .B2(net156),
    .A2(_0305_),
    .A1(_1274_));
 sg13g2_o21ai_1 _1984_ (.B1(_1274_),
    .Y(_0308_),
    .A1(net156),
    .A2(_0304_));
 sg13g2_nor2b_1 _1985_ (.A(_0306_),
    .B_N(_0308_),
    .Y(_0309_));
 sg13g2_or2_1 _1986_ (.X(_0310_),
    .B(_0309_),
    .A(net156));
 sg13g2_xnor2_1 _1987_ (.Y(_0311_),
    .A(\u_cnt0.count[4] ),
    .B(_0309_));
 sg13g2_nor2_1 _1988_ (.A(\u_cnt0.count[3] ),
    .B(_0311_),
    .Y(_0312_));
 sg13g2_a22oi_1 _1989_ (.Y(_0313_),
    .B1(_0310_),
    .B2(_0304_),
    .A2(_0306_),
    .A1(_0952_));
 sg13g2_o21ai_1 _1990_ (.B1(_0307_),
    .Y(_0314_),
    .A1(_0312_),
    .A2(_0313_));
 sg13g2_xor2_1 _1991_ (.B(_0314_),
    .A(net874),
    .X(_0315_));
 sg13g2_and2_1 _1992_ (.A(net646),
    .B(_0315_),
    .X(_0316_));
 sg13g2_o21ai_1 _1993_ (.B1(_0316_),
    .Y(_0317_),
    .A1(_1270_),
    .A2(_1271_));
 sg13g2_nand2_1 _1994_ (.Y(_0270_),
    .A(_1268_),
    .B(_0317_));
 sg13g2_xnor2_1 _1995_ (.Y(_0292_),
    .A(_0949_),
    .B(_0288_));
 sg13g2_a21oi_1 _1996_ (.A1(_0949_),
    .A2(_0288_),
    .Y(_0318_),
    .B1(_1029_));
 sg13g2_a21o_1 _1997_ (.A2(_1061_),
    .A1(_1030_),
    .B1(_0318_),
    .X(_0293_));
 sg13g2_mux2_1 _1998_ (.A0(_1061_),
    .A1(_1031_),
    .S(_1030_),
    .X(_0294_));
 sg13g2_nor2_1 _1999_ (.A(net646),
    .B(_1268_),
    .Y(_0319_));
 sg13g2_xnor2_1 _2000_ (.Y(_0274_),
    .A(_0954_),
    .B(_0270_));
 sg13g2_nand3_1 _2001_ (.B(_1269_),
    .C(_1272_),
    .A(_0954_),
    .Y(_0320_));
 sg13g2_o21ai_1 _2002_ (.B1(_0320_),
    .Y(_0275_),
    .A1(_1272_),
    .A2(_0319_));
 sg13g2_a22oi_1 _2003_ (.Y(_0321_),
    .B1(_0317_),
    .B2(_1268_),
    .A2(_1272_),
    .A1(_0954_));
 sg13g2_nand4_1 _2004_ (.B(_0307_),
    .C(_0311_),
    .A(\u_cnt0.count[3] ),
    .Y(_0322_),
    .D(_0313_));
 sg13g2_nand2b_1 _2005_ (.Y(_0323_),
    .B(_0312_),
    .A_N(_0313_));
 sg13g2_nand3_1 _2006_ (.B(_0322_),
    .C(_0323_),
    .A(_0307_),
    .Y(_0324_));
 sg13g2_and2_1 _2007_ (.A(_0953_),
    .B(_0324_),
    .X(_0325_));
 sg13g2_xnor2_1 _2008_ (.Y(_0326_),
    .A(_0315_),
    .B(_0325_));
 sg13g2_xnor2_1 _2009_ (.Y(_0276_),
    .A(_0321_),
    .B(_0326_));
 sg13g2_xnor2_1 _2010_ (.Y(_0301_),
    .A(net587),
    .B(_1128_));
 sg13g2_o21ai_1 _2011_ (.B1(_1126_),
    .Y(_0327_),
    .A1(net587),
    .A2(_1128_));
 sg13g2_nor2_1 _2012_ (.A(net587),
    .B(_1126_),
    .Y(_0328_));
 sg13g2_nand2_1 _2013_ (.Y(_0329_),
    .A(_1125_),
    .B(_0328_));
 sg13g2_nand2_1 _2014_ (.Y(_0302_),
    .A(_0327_),
    .B(_0329_));
 sg13g2_nor2_1 _2015_ (.A(_1128_),
    .B(_0328_),
    .Y(_0330_));
 sg13g2_xnor2_1 _2016_ (.Y(_0331_),
    .A(_1115_),
    .B(_1124_));
 sg13g2_xnor2_1 _2017_ (.Y(_0303_),
    .A(_0330_),
    .B(_0331_));
 sg13g2_nor2_1 _2018_ (.A(net595),
    .B(_1198_),
    .Y(_0332_));
 sg13g2_xnor2_1 _2019_ (.Y(_0283_),
    .A(net595),
    .B(_1198_));
 sg13g2_xor2_1 _2020_ (.B(_0332_),
    .A(_1193_),
    .X(_0284_));
 sg13g2_o21ai_1 _2021_ (.B1(_0279_),
    .Y(_0333_),
    .A1(net595),
    .A2(_1193_));
 sg13g2_nand3b_1 _2022_ (.B(_1186_),
    .C(_0951_),
    .Y(_0334_),
    .A_N(_1184_));
 sg13g2_nand2_1 _2023_ (.Y(_0335_),
    .A(_1192_),
    .B(_0334_));
 sg13g2_xnor2_1 _2024_ (.Y(_0285_),
    .A(_0333_),
    .B(_0335_));
 sg13g2_and2_1 _2025_ (.A(net561),
    .B(_0981_),
    .X(_0001_));
 sg13g2_and4_1 _2026_ (.A(net606),
    .B(net157),
    .C(\u_uart.state[1] ),
    .D(_1079_),
    .X(_0000_));
 sg13g2_nand3_1 _2027_ (.B(\u_deb0.counter[2] ),
    .C(\u_deb0.counter[1] ),
    .A(\u_deb0.counter[3] ),
    .Y(_0336_));
 sg13g2_nand3_1 _2028_ (.B(net520),
    .C(net702),
    .A(net543),
    .Y(_0337_));
 sg13g2_nor2_1 _2029_ (.A(\u_deb0.counter[8] ),
    .B(\u_deb0.counter[7] ),
    .Y(_0338_));
 sg13g2_o21ai_1 _2030_ (.B1(_0338_),
    .Y(_0339_),
    .A1(_0336_),
    .A2(_0337_));
 sg13g2_a21oi_1 _2031_ (.A1(\u_deb0.counter[9] ),
    .A2(_0339_),
    .Y(_0340_),
    .B1(\u_deb0.counter[10] ));
 sg13g2_nand2_1 _2032_ (.Y(_0341_),
    .A(\u_deb0.counter[12] ),
    .B(\u_deb0.counter[11] ));
 sg13g2_nor4_1 _2033_ (.A(\u_deb0.counter[16] ),
    .B(\u_deb0.counter[15] ),
    .C(\u_deb0.counter[14] ),
    .D(\u_deb0.counter[13] ),
    .Y(_0342_));
 sg13g2_o21ai_1 _2034_ (.B1(_0342_),
    .Y(_0343_),
    .A1(_0340_),
    .A2(_0341_));
 sg13g2_and2_1 _2035_ (.A(net509),
    .B(net552),
    .X(_0344_));
 sg13g2_a21oi_2 _2036_ (.B1(net732),
    .Y(_0345_),
    .A2(_0344_),
    .A1(_0343_));
 sg13g2_xor2_1 _2037_ (.B(net5),
    .A(\u_deb0.Output ),
    .X(_0346_));
 sg13g2_nand3_1 _2038_ (.B(_0345_),
    .C(_0346_),
    .A(net158),
    .Y(_0347_));
 sg13g2_inv_2 _2039_ (.Y(_0348_),
    .A(net137));
 sg13g2_nor2_1 _2040_ (.A(net445),
    .B(net136),
    .Y(_0009_));
 sg13g2_xnor2_1 _2041_ (.Y(_0349_),
    .A(net743),
    .B(net445));
 sg13g2_nor2_1 _2042_ (.A(net136),
    .B(_0349_),
    .Y(_0010_));
 sg13g2_a21oi_1 _2043_ (.A1(\u_deb0.counter[1] ),
    .A2(net445),
    .Y(_0350_),
    .B1(net584));
 sg13g2_and3_1 _2044_ (.X(_0351_),
    .A(net584),
    .B(net909),
    .C(net445));
 sg13g2_nor3_1 _2045_ (.A(net136),
    .B(net585),
    .C(_0351_),
    .Y(_0011_));
 sg13g2_and2_1 _2046_ (.A(net634),
    .B(_0351_),
    .X(_0352_));
 sg13g2_nor2_1 _2047_ (.A(net634),
    .B(_0351_),
    .Y(_0353_));
 sg13g2_nor3_1 _2048_ (.A(net136),
    .B(_0352_),
    .C(net635),
    .Y(_0012_));
 sg13g2_nor2_1 _2049_ (.A(net702),
    .B(_0352_),
    .Y(_0354_));
 sg13g2_and2_1 _2050_ (.A(net702),
    .B(_0352_),
    .X(_0355_));
 sg13g2_nor3_1 _2051_ (.A(net136),
    .B(_0354_),
    .C(_0355_),
    .Y(_0013_));
 sg13g2_o21ai_1 _2052_ (.B1(_0348_),
    .Y(_0356_),
    .A1(net520),
    .A2(_0355_));
 sg13g2_a21oi_1 _2053_ (.A1(net520),
    .A2(_0355_),
    .Y(_0014_),
    .B1(_0356_));
 sg13g2_a21oi_1 _2054_ (.A1(net520),
    .A2(_0355_),
    .Y(_0357_),
    .B1(net543));
 sg13g2_nor2b_1 _2055_ (.A(_0337_),
    .B_N(_0352_),
    .Y(_0358_));
 sg13g2_nor3_1 _2056_ (.A(net136),
    .B(net544),
    .C(_0358_),
    .Y(_0015_));
 sg13g2_and2_1 _2057_ (.A(net656),
    .B(_0358_),
    .X(_0359_));
 sg13g2_nor2_1 _2058_ (.A(net656),
    .B(_0358_),
    .Y(_0360_));
 sg13g2_nor3_1 _2059_ (.A(net136),
    .B(_0359_),
    .C(net657),
    .Y(_0016_));
 sg13g2_nor2_1 _2060_ (.A(net725),
    .B(_0359_),
    .Y(_0361_));
 sg13g2_and2_1 _2061_ (.A(net725),
    .B(_0359_),
    .X(_0362_));
 sg13g2_nor3_1 _2062_ (.A(net137),
    .B(_0361_),
    .C(_0362_),
    .Y(_0017_));
 sg13g2_nor2_1 _2063_ (.A(net742),
    .B(_0362_),
    .Y(_0363_));
 sg13g2_and2_1 _2064_ (.A(net742),
    .B(_0362_),
    .X(_0364_));
 sg13g2_nor3_1 _2065_ (.A(net136),
    .B(_0363_),
    .C(_0364_),
    .Y(_0018_));
 sg13g2_and2_1 _2066_ (.A(net603),
    .B(_0364_),
    .X(_0365_));
 sg13g2_nor2_1 _2067_ (.A(net603),
    .B(_0364_),
    .Y(_0366_));
 sg13g2_nor3_1 _2068_ (.A(net137),
    .B(_0365_),
    .C(net604),
    .Y(_0019_));
 sg13g2_xnor2_1 _2069_ (.Y(_0367_),
    .A(net784),
    .B(_0365_));
 sg13g2_nor2_1 _2070_ (.A(net137),
    .B(_0367_),
    .Y(_0020_));
 sg13g2_a21oi_1 _2071_ (.A1(\u_deb0.counter[11] ),
    .A2(_0365_),
    .Y(_0368_),
    .B1(net643));
 sg13g2_and3_1 _2072_ (.X(_0369_),
    .A(net643),
    .B(net784),
    .C(_0365_));
 sg13g2_nor3_1 _2073_ (.A(net137),
    .B(net644),
    .C(_0369_),
    .Y(_0021_));
 sg13g2_and4_1 _2074_ (.A(net814),
    .B(net643),
    .C(net784),
    .D(_0365_),
    .X(_0370_));
 sg13g2_o21ai_1 _2075_ (.B1(_0348_),
    .Y(_0371_),
    .A1(net814),
    .A2(_0369_));
 sg13g2_nor2_1 _2076_ (.A(_0370_),
    .B(_0371_),
    .Y(_0022_));
 sg13g2_and2_1 _2077_ (.A(net844),
    .B(_0370_),
    .X(_0372_));
 sg13g2_o21ai_1 _2078_ (.B1(_0348_),
    .Y(_0373_),
    .A1(net844),
    .A2(_0370_));
 sg13g2_nor2_1 _2079_ (.A(_0372_),
    .B(_0373_),
    .Y(_0023_));
 sg13g2_and2_1 _2080_ (.A(net821),
    .B(_0372_),
    .X(_0374_));
 sg13g2_o21ai_1 _2081_ (.B1(_0348_),
    .Y(_0375_),
    .A1(net821),
    .A2(_0372_));
 sg13g2_nor2_1 _2082_ (.A(_0374_),
    .B(net822),
    .Y(_0024_));
 sg13g2_nor2_1 _2083_ (.A(net676),
    .B(_0374_),
    .Y(_0376_));
 sg13g2_and2_1 _2084_ (.A(net676),
    .B(_0374_),
    .X(_0377_));
 sg13g2_nor3_1 _2085_ (.A(net137),
    .B(net677),
    .C(_0377_),
    .Y(_0025_));
 sg13g2_o21ai_1 _2086_ (.B1(_0348_),
    .Y(_0378_),
    .A1(net552),
    .A2(_0377_));
 sg13g2_a21oi_1 _2087_ (.A1(net552),
    .A2(_0377_),
    .Y(_0026_),
    .B1(_0378_));
 sg13g2_a21oi_1 _2088_ (.A1(\u_deb0.counter[17] ),
    .A2(_0377_),
    .Y(_0379_),
    .B1(net509));
 sg13g2_nor2_1 _2089_ (.A(net137),
    .B(net510),
    .Y(_0027_));
 sg13g2_o21ai_1 _2090_ (.B1(net159),
    .Y(_0380_),
    .A1(net5),
    .A2(_0345_));
 sg13g2_a21oi_1 _2091_ (.A1(_0959_),
    .A2(net733),
    .Y(_0029_),
    .B1(_0380_));
 sg13g2_nand3_1 _2092_ (.B(\u_deb1.counter[2] ),
    .C(\u_deb1.counter[1] ),
    .A(\u_deb1.counter[3] ),
    .Y(_0381_));
 sg13g2_nand3_1 _2093_ (.B(net513),
    .C(\u_deb1.counter[4] ),
    .A(net538),
    .Y(_0382_));
 sg13g2_nor2_1 _2094_ (.A(\u_deb1.counter[8] ),
    .B(\u_deb1.counter[7] ),
    .Y(_0383_));
 sg13g2_o21ai_1 _2095_ (.B1(_0383_),
    .Y(_0384_),
    .A1(_0381_),
    .A2(_0382_));
 sg13g2_a21oi_1 _2096_ (.A1(\u_deb1.counter[9] ),
    .A2(_0384_),
    .Y(_0385_),
    .B1(net682));
 sg13g2_nand2_1 _2097_ (.Y(_0386_),
    .A(net628),
    .B(net788));
 sg13g2_nor4_1 _2098_ (.A(net753),
    .B(net834),
    .C(net806),
    .D(net835),
    .Y(_0387_));
 sg13g2_o21ai_1 _2099_ (.B1(_0387_),
    .Y(_0388_),
    .A1(_0385_),
    .A2(_0386_));
 sg13g2_and2_1 _2100_ (.A(net524),
    .B(net546),
    .X(_0389_));
 sg13g2_a21oi_1 _2101_ (.A1(_0388_),
    .A2(_0389_),
    .Y(_0390_),
    .B1(net839));
 sg13g2_xor2_1 _2102_ (.B(net1),
    .A(net765),
    .X(_0391_));
 sg13g2_nand3_1 _2103_ (.B(_0390_),
    .C(_0391_),
    .A(net159),
    .Y(_0392_));
 sg13g2_inv_2 _2104_ (.Y(_0393_),
    .A(net134));
 sg13g2_nor2_1 _2105_ (.A(net463),
    .B(net135),
    .Y(_0030_));
 sg13g2_xnor2_1 _2106_ (.Y(_0394_),
    .A(net712),
    .B(net463));
 sg13g2_nor2_1 _2107_ (.A(net134),
    .B(_0394_),
    .Y(_0031_));
 sg13g2_a21oi_1 _2108_ (.A1(\u_deb1.counter[1] ),
    .A2(net463),
    .Y(_0395_),
    .B1(net580));
 sg13g2_and3_1 _2109_ (.X(_0396_),
    .A(net580),
    .B(\u_deb1.counter[1] ),
    .C(net463));
 sg13g2_nor3_1 _2110_ (.A(net135),
    .B(net581),
    .C(_0396_),
    .Y(_0032_));
 sg13g2_and2_1 _2111_ (.A(net619),
    .B(_0396_),
    .X(_0397_));
 sg13g2_nor2_1 _2112_ (.A(net619),
    .B(_0396_),
    .Y(_0398_));
 sg13g2_nor3_1 _2113_ (.A(net135),
    .B(_0397_),
    .C(net620),
    .Y(_0033_));
 sg13g2_nor2_1 _2114_ (.A(net710),
    .B(_0397_),
    .Y(_0399_));
 sg13g2_and2_1 _2115_ (.A(net710),
    .B(_0397_),
    .X(_0400_));
 sg13g2_nor3_1 _2116_ (.A(net135),
    .B(_0399_),
    .C(_0400_),
    .Y(_0034_));
 sg13g2_o21ai_1 _2117_ (.B1(_0393_),
    .Y(_0401_),
    .A1(net513),
    .A2(_0400_));
 sg13g2_a21oi_1 _2118_ (.A1(net513),
    .A2(_0400_),
    .Y(_0035_),
    .B1(_0401_));
 sg13g2_a21oi_1 _2119_ (.A1(net513),
    .A2(_0400_),
    .Y(_0402_),
    .B1(net538));
 sg13g2_nor2b_1 _2120_ (.A(_0382_),
    .B_N(_0397_),
    .Y(_0403_));
 sg13g2_nor3_1 _2121_ (.A(net135),
    .B(net539),
    .C(_0403_),
    .Y(_0036_));
 sg13g2_and2_1 _2122_ (.A(net616),
    .B(_0403_),
    .X(_0404_));
 sg13g2_nor2_1 _2123_ (.A(net616),
    .B(_0403_),
    .Y(_0405_));
 sg13g2_nor3_1 _2124_ (.A(net135),
    .B(_0404_),
    .C(net617),
    .Y(_0037_));
 sg13g2_nor2_1 _2125_ (.A(net692),
    .B(_0404_),
    .Y(_0406_));
 sg13g2_and2_1 _2126_ (.A(net692),
    .B(_0404_),
    .X(_0407_));
 sg13g2_nor3_1 _2127_ (.A(net135),
    .B(net693),
    .C(_0407_),
    .Y(_0038_));
 sg13g2_nor2_1 _2128_ (.A(net697),
    .B(_0407_),
    .Y(_0408_));
 sg13g2_and2_1 _2129_ (.A(net697),
    .B(_0407_),
    .X(_0409_));
 sg13g2_nor3_1 _2130_ (.A(net134),
    .B(_0408_),
    .C(_0409_),
    .Y(_0039_));
 sg13g2_and2_1 _2131_ (.A(net682),
    .B(_0409_),
    .X(_0410_));
 sg13g2_nor2_1 _2132_ (.A(net682),
    .B(_0409_),
    .Y(_0411_));
 sg13g2_nor3_1 _2133_ (.A(net134),
    .B(_0410_),
    .C(net683),
    .Y(_0040_));
 sg13g2_xnor2_1 _2134_ (.Y(_0412_),
    .A(net788),
    .B(_0410_));
 sg13g2_nor2_1 _2135_ (.A(net134),
    .B(_0412_),
    .Y(_0041_));
 sg13g2_a21oi_1 _2136_ (.A1(\u_deb1.counter[11] ),
    .A2(_0410_),
    .Y(_0413_),
    .B1(net628));
 sg13g2_and3_1 _2137_ (.X(_0414_),
    .A(net628),
    .B(net788),
    .C(_0410_));
 sg13g2_nor3_1 _2138_ (.A(net134),
    .B(net629),
    .C(_0414_),
    .Y(_0042_));
 sg13g2_and4_1 _2139_ (.A(net835),
    .B(net628),
    .C(net788),
    .D(_0410_),
    .X(_0415_));
 sg13g2_o21ai_1 _2140_ (.B1(_0393_),
    .Y(_0416_),
    .A1(net835),
    .A2(_0414_));
 sg13g2_nor2_1 _2141_ (.A(_0415_),
    .B(_0416_),
    .Y(_0043_));
 sg13g2_and2_1 _2142_ (.A(net806),
    .B(_0415_),
    .X(_0417_));
 sg13g2_o21ai_1 _2143_ (.B1(_0393_),
    .Y(_0418_),
    .A1(net806),
    .A2(_0415_));
 sg13g2_nor2_1 _2144_ (.A(_0417_),
    .B(net807),
    .Y(_0044_));
 sg13g2_and2_1 _2145_ (.A(net834),
    .B(_0417_),
    .X(_0419_));
 sg13g2_o21ai_1 _2146_ (.B1(_0393_),
    .Y(_0420_),
    .A1(net834),
    .A2(_0417_));
 sg13g2_nor2_1 _2147_ (.A(_0419_),
    .B(_0420_),
    .Y(_0045_));
 sg13g2_nor2_1 _2148_ (.A(net753),
    .B(_0419_),
    .Y(_0421_));
 sg13g2_and2_1 _2149_ (.A(net753),
    .B(_0419_),
    .X(_0422_));
 sg13g2_nor3_1 _2150_ (.A(net134),
    .B(net754),
    .C(_0422_),
    .Y(_0046_));
 sg13g2_o21ai_1 _2151_ (.B1(_0393_),
    .Y(_0423_),
    .A1(net546),
    .A2(_0422_));
 sg13g2_a21oi_1 _2152_ (.A1(net546),
    .A2(_0422_),
    .Y(_0047_),
    .B1(_0423_));
 sg13g2_a21oi_1 _2153_ (.A1(\u_deb1.counter[17] ),
    .A2(_0422_),
    .Y(_0424_),
    .B1(net524));
 sg13g2_nor2_1 _2154_ (.A(net134),
    .B(net525),
    .Y(_0048_));
 sg13g2_o21ai_1 _2155_ (.B1(net159),
    .Y(_0425_),
    .A1(net1),
    .A2(_0390_));
 sg13g2_a21oi_1 _2156_ (.A1(_0958_),
    .A2(_0390_),
    .Y(_0050_),
    .B1(_0425_));
 sg13g2_nand3_1 _2157_ (.B(\u_deb2.counter[2] ),
    .C(\u_deb2.counter[1] ),
    .A(\u_deb2.counter[3] ),
    .Y(_0426_));
 sg13g2_nand3_1 _2158_ (.B(net515),
    .C(\u_deb2.counter[4] ),
    .A(net558),
    .Y(_0427_));
 sg13g2_nor2_1 _2159_ (.A(\u_deb2.counter[8] ),
    .B(\u_deb2.counter[7] ),
    .Y(_0428_));
 sg13g2_o21ai_1 _2160_ (.B1(_0428_),
    .Y(_0429_),
    .A1(_0426_),
    .A2(_0427_));
 sg13g2_a21oi_1 _2161_ (.A1(\u_deb2.counter[9] ),
    .A2(_0429_),
    .Y(_0430_),
    .B1(\u_deb2.counter[10] ));
 sg13g2_nand2_1 _2162_ (.Y(_0431_),
    .A(net600),
    .B(\u_deb2.counter[11] ));
 sg13g2_nor4_1 _2163_ (.A(\u_deb2.counter[16] ),
    .B(\u_deb2.counter[15] ),
    .C(\u_deb2.counter[14] ),
    .D(\u_deb2.counter[13] ),
    .Y(_0432_));
 sg13g2_o21ai_1 _2164_ (.B1(_0432_),
    .Y(_0433_),
    .A1(_0430_),
    .A2(_0431_));
 sg13g2_and2_1 _2165_ (.A(net527),
    .B(net556),
    .X(_0434_));
 sg13g2_a21oi_1 _2166_ (.A1(_0433_),
    .A2(_0434_),
    .Y(_0435_),
    .B1(net695));
 sg13g2_xor2_1 _2167_ (.B(net2),
    .A(net573),
    .X(_0436_));
 sg13g2_nand3_1 _2168_ (.B(_0435_),
    .C(_0436_),
    .A(net159),
    .Y(_0437_));
 sg13g2_inv_2 _2169_ (.Y(_0438_),
    .A(net132));
 sg13g2_nor2_1 _2170_ (.A(net469),
    .B(net133),
    .Y(_0051_));
 sg13g2_xnor2_1 _2171_ (.Y(_0439_),
    .A(net731),
    .B(net469));
 sg13g2_nor2_1 _2172_ (.A(net133),
    .B(_0439_),
    .Y(_0052_));
 sg13g2_a21oi_1 _2173_ (.A1(\u_deb2.counter[1] ),
    .A2(net469),
    .Y(_0440_),
    .B1(net574));
 sg13g2_and3_1 _2174_ (.X(_0441_),
    .A(net574),
    .B(net908),
    .C(net469));
 sg13g2_nor3_1 _2175_ (.A(net132),
    .B(net575),
    .C(_0441_),
    .Y(_0053_));
 sg13g2_and2_1 _2176_ (.A(net653),
    .B(_0441_),
    .X(_0442_));
 sg13g2_nor2_1 _2177_ (.A(net653),
    .B(_0441_),
    .Y(_0443_));
 sg13g2_nor3_1 _2178_ (.A(net133),
    .B(_0442_),
    .C(net654),
    .Y(_0054_));
 sg13g2_nor2_1 _2179_ (.A(net727),
    .B(_0442_),
    .Y(_0444_));
 sg13g2_and2_1 _2180_ (.A(net727),
    .B(_0442_),
    .X(_0445_));
 sg13g2_nor3_1 _2181_ (.A(net133),
    .B(_0444_),
    .C(_0445_),
    .Y(_0055_));
 sg13g2_o21ai_1 _2182_ (.B1(_0438_),
    .Y(_0446_),
    .A1(net515),
    .A2(_0445_));
 sg13g2_a21oi_1 _2183_ (.A1(net515),
    .A2(_0445_),
    .Y(_0056_),
    .B1(_0446_));
 sg13g2_a21oi_1 _2184_ (.A1(net515),
    .A2(_0445_),
    .Y(_0447_),
    .B1(net558));
 sg13g2_nor2b_1 _2185_ (.A(_0427_),
    .B_N(_0442_),
    .Y(_0448_));
 sg13g2_nor3_1 _2186_ (.A(net133),
    .B(net559),
    .C(_0448_),
    .Y(_0057_));
 sg13g2_and2_1 _2187_ (.A(net650),
    .B(_0448_),
    .X(_0449_));
 sg13g2_nor2_1 _2188_ (.A(net650),
    .B(_0448_),
    .Y(_0450_));
 sg13g2_nor3_1 _2189_ (.A(net133),
    .B(_0449_),
    .C(net651),
    .Y(_0058_));
 sg13g2_nor2_1 _2190_ (.A(net689),
    .B(_0449_),
    .Y(_0451_));
 sg13g2_and2_1 _2191_ (.A(net689),
    .B(_0449_),
    .X(_0452_));
 sg13g2_nor3_1 _2192_ (.A(net133),
    .B(net690),
    .C(_0452_),
    .Y(_0059_));
 sg13g2_nor2_1 _2193_ (.A(net709),
    .B(_0452_),
    .Y(_0453_));
 sg13g2_and2_1 _2194_ (.A(net709),
    .B(_0452_),
    .X(_0454_));
 sg13g2_nor3_1 _2195_ (.A(net132),
    .B(_0453_),
    .C(_0454_),
    .Y(_0060_));
 sg13g2_and2_1 _2196_ (.A(net658),
    .B(_0454_),
    .X(_0455_));
 sg13g2_nor2_1 _2197_ (.A(net658),
    .B(_0454_),
    .Y(_0456_));
 sg13g2_nor3_1 _2198_ (.A(net132),
    .B(_0455_),
    .C(net659),
    .Y(_0061_));
 sg13g2_xnor2_1 _2199_ (.Y(_0457_),
    .A(net798),
    .B(_0455_));
 sg13g2_nor2_1 _2200_ (.A(net132),
    .B(_0457_),
    .Y(_0062_));
 sg13g2_a21oi_1 _2201_ (.A1(\u_deb2.counter[11] ),
    .A2(_0455_),
    .Y(_0458_),
    .B1(net600));
 sg13g2_and3_1 _2202_ (.X(_0459_),
    .A(net600),
    .B(net798),
    .C(_0455_));
 sg13g2_nor3_1 _2203_ (.A(net132),
    .B(net601),
    .C(_0459_),
    .Y(_0063_));
 sg13g2_and4_1 _2204_ (.A(net817),
    .B(net600),
    .C(net798),
    .D(_0455_),
    .X(_0460_));
 sg13g2_o21ai_1 _2205_ (.B1(_0438_),
    .Y(_0461_),
    .A1(net817),
    .A2(_0459_));
 sg13g2_nor2_1 _2206_ (.A(_0460_),
    .B(_0461_),
    .Y(_0064_));
 sg13g2_and2_1 _2207_ (.A(net818),
    .B(_0460_),
    .X(_0462_));
 sg13g2_o21ai_1 _2208_ (.B1(_0438_),
    .Y(_0463_),
    .A1(net818),
    .A2(_0460_));
 sg13g2_nor2_1 _2209_ (.A(_0462_),
    .B(_0463_),
    .Y(_0065_));
 sg13g2_and2_1 _2210_ (.A(net838),
    .B(_0462_),
    .X(_0464_));
 sg13g2_o21ai_1 _2211_ (.B1(_0438_),
    .Y(_0465_),
    .A1(net838),
    .A2(_0462_));
 sg13g2_nor2_1 _2212_ (.A(_0464_),
    .B(_0465_),
    .Y(_0066_));
 sg13g2_nor2_1 _2213_ (.A(net737),
    .B(_0464_),
    .Y(_0466_));
 sg13g2_and2_1 _2214_ (.A(net737),
    .B(_0464_),
    .X(_0467_));
 sg13g2_nor3_1 _2215_ (.A(net132),
    .B(net738),
    .C(_0467_),
    .Y(_0067_));
 sg13g2_o21ai_1 _2216_ (.B1(_0438_),
    .Y(_0468_),
    .A1(net556),
    .A2(_0467_));
 sg13g2_a21oi_1 _2217_ (.A1(net556),
    .A2(_0467_),
    .Y(_0068_),
    .B1(_0468_));
 sg13g2_a21oi_1 _2218_ (.A1(\u_deb2.counter[17] ),
    .A2(_0467_),
    .Y(_0469_),
    .B1(net527));
 sg13g2_nor2_1 _2219_ (.A(net132),
    .B(net528),
    .Y(_0069_));
 sg13g2_o21ai_1 _2220_ (.B1(net159),
    .Y(_0470_),
    .A1(net2),
    .A2(net696));
 sg13g2_a21oi_1 _2221_ (.A1(_0957_),
    .A2(net696),
    .Y(_0071_),
    .B1(_0470_));
 sg13g2_nand3_1 _2222_ (.B(\u_deb3.counter[2] ),
    .C(\u_deb3.counter[1] ),
    .A(\u_deb3.counter[3] ),
    .Y(_0471_));
 sg13g2_nand3_1 _2223_ (.B(net522),
    .C(net904),
    .A(net530),
    .Y(_0472_));
 sg13g2_nor2_1 _2224_ (.A(\u_deb3.counter[8] ),
    .B(\u_deb3.counter[7] ),
    .Y(_0473_));
 sg13g2_o21ai_1 _2225_ (.B1(_0473_),
    .Y(_0474_),
    .A1(_0471_),
    .A2(_0472_));
 sg13g2_a21oi_1 _2226_ (.A1(\u_deb3.counter[9] ),
    .A2(_0474_),
    .Y(_0475_),
    .B1(net706));
 sg13g2_nand2_1 _2227_ (.Y(_0476_),
    .A(net608),
    .B(\u_deb3.counter[11] ));
 sg13g2_nor4_1 _2228_ (.A(net699),
    .B(\u_deb3.counter[15] ),
    .C(\u_deb3.counter[14] ),
    .D(\u_deb3.counter[13] ),
    .Y(_0477_));
 sg13g2_o21ai_1 _2229_ (.B1(_0477_),
    .Y(_0478_),
    .A1(_0475_),
    .A2(_0476_));
 sg13g2_and2_1 _2230_ (.A(net517),
    .B(net550),
    .X(_0479_));
 sg13g2_a21oi_1 _2231_ (.A1(_0478_),
    .A2(_0479_),
    .Y(_0480_),
    .B1(net720));
 sg13g2_xor2_1 _2232_ (.B(net3),
    .A(net583),
    .X(_0481_));
 sg13g2_nand3_1 _2233_ (.B(_0480_),
    .C(_0481_),
    .A(net159),
    .Y(_0482_));
 sg13g2_inv_2 _2234_ (.Y(_0483_),
    .A(net130));
 sg13g2_nor2_1 _2235_ (.A(net456),
    .B(net130),
    .Y(_0072_));
 sg13g2_xnor2_1 _2236_ (.Y(_0484_),
    .A(net740),
    .B(net456));
 sg13g2_nor2_1 _2237_ (.A(net130),
    .B(_0484_),
    .Y(_0073_));
 sg13g2_a21oi_1 _2238_ (.A1(\u_deb3.counter[1] ),
    .A2(net456),
    .Y(_0485_),
    .B1(net568));
 sg13g2_and3_1 _2239_ (.X(_0486_),
    .A(net568),
    .B(\u_deb3.counter[1] ),
    .C(net456));
 sg13g2_nor3_1 _2240_ (.A(net130),
    .B(net569),
    .C(_0486_),
    .Y(_0074_));
 sg13g2_and2_1 _2241_ (.A(net622),
    .B(_0486_),
    .X(_0487_));
 sg13g2_nor2_1 _2242_ (.A(net622),
    .B(_0486_),
    .Y(_0488_));
 sg13g2_nor3_1 _2243_ (.A(net130),
    .B(_0487_),
    .C(net623),
    .Y(_0075_));
 sg13g2_nor2_1 _2244_ (.A(net764),
    .B(_0487_),
    .Y(_0489_));
 sg13g2_and2_1 _2245_ (.A(net764),
    .B(_0487_),
    .X(_0490_));
 sg13g2_nor3_1 _2246_ (.A(net131),
    .B(_0489_),
    .C(_0490_),
    .Y(_0076_));
 sg13g2_o21ai_1 _2247_ (.B1(_0483_),
    .Y(_0491_),
    .A1(net522),
    .A2(_0490_));
 sg13g2_a21oi_1 _2248_ (.A1(net522),
    .A2(_0490_),
    .Y(_0077_),
    .B1(_0491_));
 sg13g2_a21oi_1 _2249_ (.A1(net522),
    .A2(_0490_),
    .Y(_0492_),
    .B1(net530));
 sg13g2_nor2b_1 _2250_ (.A(_0472_),
    .B_N(_0487_),
    .Y(_0493_));
 sg13g2_nor3_1 _2251_ (.A(net131),
    .B(net531),
    .C(_0493_),
    .Y(_0078_));
 sg13g2_and2_1 _2252_ (.A(net679),
    .B(_0493_),
    .X(_0494_));
 sg13g2_nor2_1 _2253_ (.A(net679),
    .B(_0493_),
    .Y(_0495_));
 sg13g2_nor3_1 _2254_ (.A(net131),
    .B(_0494_),
    .C(net680),
    .Y(_0079_));
 sg13g2_nor2_1 _2255_ (.A(net741),
    .B(_0494_),
    .Y(_0496_));
 sg13g2_and2_1 _2256_ (.A(net741),
    .B(_0494_),
    .X(_0497_));
 sg13g2_nor3_1 _2257_ (.A(net131),
    .B(_0496_),
    .C(_0497_),
    .Y(_0080_));
 sg13g2_nor2_1 _2258_ (.A(net664),
    .B(_0497_),
    .Y(_0498_));
 sg13g2_and2_1 _2259_ (.A(net664),
    .B(_0497_),
    .X(_0499_));
 sg13g2_nor3_1 _2260_ (.A(net131),
    .B(net665),
    .C(_0499_),
    .Y(_0081_));
 sg13g2_and2_1 _2261_ (.A(net706),
    .B(_0499_),
    .X(_0500_));
 sg13g2_nor2_1 _2262_ (.A(net706),
    .B(_0499_),
    .Y(_0501_));
 sg13g2_nor3_1 _2263_ (.A(net130),
    .B(_0500_),
    .C(net707),
    .Y(_0082_));
 sg13g2_xnor2_1 _2264_ (.Y(_0502_),
    .A(net819),
    .B(_0500_));
 sg13g2_nor2_1 _2265_ (.A(net131),
    .B(_0502_),
    .Y(_0083_));
 sg13g2_a21oi_1 _2266_ (.A1(\u_deb3.counter[11] ),
    .A2(_0500_),
    .Y(_0503_),
    .B1(net608));
 sg13g2_and3_1 _2267_ (.X(_0504_),
    .A(net608),
    .B(net819),
    .C(_0500_));
 sg13g2_nor3_1 _2268_ (.A(net131),
    .B(net609),
    .C(_0504_),
    .Y(_0084_));
 sg13g2_and4_1 _2269_ (.A(net845),
    .B(net608),
    .C(net819),
    .D(_0500_),
    .X(_0505_));
 sg13g2_o21ai_1 _2270_ (.B1(_0483_),
    .Y(_0506_),
    .A1(net845),
    .A2(_0504_));
 sg13g2_nor2_1 _2271_ (.A(_0505_),
    .B(_0506_),
    .Y(_0085_));
 sg13g2_and2_1 _2272_ (.A(net811),
    .B(_0505_),
    .X(_0507_));
 sg13g2_o21ai_1 _2273_ (.B1(_0483_),
    .Y(_0508_),
    .A1(net811),
    .A2(_0505_));
 sg13g2_nor2_1 _2274_ (.A(_0507_),
    .B(net812),
    .Y(_0086_));
 sg13g2_and2_1 _2275_ (.A(net830),
    .B(_0507_),
    .X(_0509_));
 sg13g2_o21ai_1 _2276_ (.B1(_0483_),
    .Y(_0510_),
    .A1(net830),
    .A2(_0507_));
 sg13g2_nor2_1 _2277_ (.A(_0509_),
    .B(_0510_),
    .Y(_0087_));
 sg13g2_nor2_1 _2278_ (.A(net699),
    .B(_0509_),
    .Y(_0511_));
 sg13g2_and2_1 _2279_ (.A(net699),
    .B(_0509_),
    .X(_0512_));
 sg13g2_nor3_1 _2280_ (.A(net130),
    .B(net700),
    .C(_0512_),
    .Y(_0088_));
 sg13g2_o21ai_1 _2281_ (.B1(_0483_),
    .Y(_0513_),
    .A1(net550),
    .A2(_0512_));
 sg13g2_a21oi_1 _2282_ (.A1(net550),
    .A2(_0512_),
    .Y(_0089_),
    .B1(_0513_));
 sg13g2_a21oi_1 _2283_ (.A1(\u_deb3.counter[17] ),
    .A2(_0512_),
    .Y(_0514_),
    .B1(net517));
 sg13g2_nor2_1 _2284_ (.A(net130),
    .B(net518),
    .Y(_0090_));
 sg13g2_o21ai_1 _2285_ (.B1(net159),
    .Y(_0515_),
    .A1(net3),
    .A2(_0480_));
 sg13g2_a21oi_1 _2286_ (.A1(_0956_),
    .A2(net721),
    .Y(_0092_),
    .B1(_0515_));
 sg13g2_nand3_1 _2287_ (.B(\u_deb4.counter[2] ),
    .C(\u_deb4.counter[1] ),
    .A(\u_deb4.counter[3] ),
    .Y(_0516_));
 sg13g2_nand3_1 _2288_ (.B(net507),
    .C(\u_deb4.counter[4] ),
    .A(net533),
    .Y(_0517_));
 sg13g2_nor2_1 _2289_ (.A(\u_deb4.counter[8] ),
    .B(\u_deb4.counter[7] ),
    .Y(_0518_));
 sg13g2_o21ai_1 _2290_ (.B1(_0518_),
    .Y(_0519_),
    .A1(_0516_),
    .A2(_0517_));
 sg13g2_a21oi_1 _2291_ (.A1(\u_deb4.counter[9] ),
    .A2(_0519_),
    .Y(_0520_),
    .B1(\u_deb4.counter[10] ));
 sg13g2_nand2_1 _2292_ (.Y(_0521_),
    .A(net647),
    .B(\u_deb4.counter[11] ));
 sg13g2_nor4_1 _2293_ (.A(net703),
    .B(\u_deb4.counter[15] ),
    .C(\u_deb4.counter[14] ),
    .D(\u_deb4.counter[13] ),
    .Y(_0522_));
 sg13g2_o21ai_1 _2294_ (.B1(_0522_),
    .Y(_0523_),
    .A1(_0520_),
    .A2(_0521_));
 sg13g2_and2_1 _2295_ (.A(net503),
    .B(net554),
    .X(_0524_));
 sg13g2_a21oi_1 _2296_ (.A1(_0523_),
    .A2(_0524_),
    .Y(_0525_),
    .B1(net746));
 sg13g2_xor2_1 _2297_ (.B(net4),
    .A(net588),
    .X(_0526_));
 sg13g2_nand3_1 _2298_ (.B(_0525_),
    .C(_0526_),
    .A(net158),
    .Y(_0527_));
 sg13g2_inv_2 _2299_ (.Y(_0528_),
    .A(net129));
 sg13g2_nor2_1 _2300_ (.A(net449),
    .B(net128),
    .Y(_0093_));
 sg13g2_xnor2_1 _2301_ (.Y(_0529_),
    .A(net685),
    .B(net449));
 sg13g2_nor2_1 _2302_ (.A(net128),
    .B(_0529_),
    .Y(_0094_));
 sg13g2_a21oi_1 _2303_ (.A1(\u_deb4.counter[1] ),
    .A2(net449),
    .Y(_0530_),
    .B1(net577));
 sg13g2_and3_1 _2304_ (.X(_0531_),
    .A(net577),
    .B(\u_deb4.counter[1] ),
    .C(net449));
 sg13g2_nor3_1 _2305_ (.A(net128),
    .B(net578),
    .C(_0531_),
    .Y(_0095_));
 sg13g2_and2_1 _2306_ (.A(net631),
    .B(_0531_),
    .X(_0532_));
 sg13g2_nor2_1 _2307_ (.A(net631),
    .B(_0531_),
    .Y(_0533_));
 sg13g2_nor3_1 _2308_ (.A(net128),
    .B(_0532_),
    .C(net632),
    .Y(_0096_));
 sg13g2_nor2_1 _2309_ (.A(net673),
    .B(_0532_),
    .Y(_0534_));
 sg13g2_and2_1 _2310_ (.A(net673),
    .B(_0532_),
    .X(_0535_));
 sg13g2_nor3_1 _2311_ (.A(net128),
    .B(net674),
    .C(_0535_),
    .Y(_0097_));
 sg13g2_o21ai_1 _2312_ (.B1(_0528_),
    .Y(_0536_),
    .A1(net507),
    .A2(_0535_));
 sg13g2_a21oi_1 _2313_ (.A1(net507),
    .A2(_0535_),
    .Y(_0098_),
    .B1(_0536_));
 sg13g2_a21oi_1 _2314_ (.A1(net507),
    .A2(_0535_),
    .Y(_0537_),
    .B1(net533));
 sg13g2_nor2b_1 _2315_ (.A(_0517_),
    .B_N(_0532_),
    .Y(_0538_));
 sg13g2_nor3_1 _2316_ (.A(net128),
    .B(net534),
    .C(_0538_),
    .Y(_0099_));
 sg13g2_and2_1 _2317_ (.A(net661),
    .B(_0538_),
    .X(_0539_));
 sg13g2_nor2_1 _2318_ (.A(net661),
    .B(_0538_),
    .Y(_0540_));
 sg13g2_nor3_1 _2319_ (.A(net129),
    .B(_0539_),
    .C(net662),
    .Y(_0100_));
 sg13g2_nor2_1 _2320_ (.A(net670),
    .B(_0539_),
    .Y(_0541_));
 sg13g2_and2_1 _2321_ (.A(net670),
    .B(_0539_),
    .X(_0542_));
 sg13g2_nor3_1 _2322_ (.A(net128),
    .B(net671),
    .C(_0542_),
    .Y(_0101_));
 sg13g2_nor2_1 _2323_ (.A(net667),
    .B(_0542_),
    .Y(_0543_));
 sg13g2_and2_1 _2324_ (.A(net667),
    .B(_0542_),
    .X(_0544_));
 sg13g2_nor3_1 _2325_ (.A(net128),
    .B(net668),
    .C(_0544_),
    .Y(_0102_));
 sg13g2_and2_1 _2326_ (.A(net625),
    .B(_0544_),
    .X(_0545_));
 sg13g2_nor2_1 _2327_ (.A(net625),
    .B(_0544_),
    .Y(_0546_));
 sg13g2_nor3_1 _2328_ (.A(net129),
    .B(_0545_),
    .C(net626),
    .Y(_0103_));
 sg13g2_xnor2_1 _2329_ (.Y(_0547_),
    .A(net797),
    .B(_0545_));
 sg13g2_nor2_1 _2330_ (.A(net129),
    .B(_0547_),
    .Y(_0104_));
 sg13g2_a21oi_1 _2331_ (.A1(\u_deb4.counter[11] ),
    .A2(_0545_),
    .Y(_0548_),
    .B1(net647));
 sg13g2_and3_1 _2332_ (.X(_0549_),
    .A(net647),
    .B(net797),
    .C(_0545_));
 sg13g2_nor3_1 _2333_ (.A(net129),
    .B(net648),
    .C(_0549_),
    .Y(_0105_));
 sg13g2_and4_1 _2334_ (.A(net840),
    .B(net647),
    .C(net797),
    .D(_0545_),
    .X(_0550_));
 sg13g2_o21ai_1 _2335_ (.B1(_0528_),
    .Y(_0551_),
    .A1(net840),
    .A2(_0549_));
 sg13g2_nor2_1 _2336_ (.A(_0550_),
    .B(_0551_),
    .Y(_0106_));
 sg13g2_and2_1 _2337_ (.A(net827),
    .B(_0550_),
    .X(_0552_));
 sg13g2_o21ai_1 _2338_ (.B1(_0528_),
    .Y(_0553_),
    .A1(net827),
    .A2(_0550_));
 sg13g2_nor2_1 _2339_ (.A(_0552_),
    .B(net828),
    .Y(_0107_));
 sg13g2_and2_1 _2340_ (.A(net841),
    .B(_0552_),
    .X(_0554_));
 sg13g2_o21ai_1 _2341_ (.B1(_0528_),
    .Y(_0555_),
    .A1(net841),
    .A2(_0552_));
 sg13g2_nor2_1 _2342_ (.A(_0554_),
    .B(_0555_),
    .Y(_0108_));
 sg13g2_nor2_1 _2343_ (.A(net703),
    .B(_0554_),
    .Y(_0556_));
 sg13g2_and2_1 _2344_ (.A(net703),
    .B(_0554_),
    .X(_0557_));
 sg13g2_nor3_1 _2345_ (.A(net129),
    .B(net704),
    .C(_0557_),
    .Y(_0109_));
 sg13g2_o21ai_1 _2346_ (.B1(_0528_),
    .Y(_0558_),
    .A1(net554),
    .A2(_0557_));
 sg13g2_a21oi_1 _2347_ (.A1(net554),
    .A2(_0557_),
    .Y(_0110_),
    .B1(_0558_));
 sg13g2_a21oi_1 _2348_ (.A1(\u_deb4.counter[17] ),
    .A2(_0557_),
    .Y(_0559_),
    .B1(net503));
 sg13g2_nor2_1 _2349_ (.A(net129),
    .B(net504),
    .Y(_0111_));
 sg13g2_o21ai_1 _2350_ (.B1(net157),
    .Y(_0560_),
    .A1(net4),
    .A2(net747));
 sg13g2_a21oi_1 _2351_ (.A1(_0955_),
    .A2(net747),
    .Y(_0113_),
    .B1(_0560_));
 sg13g2_nor2_1 _2352_ (.A(change0),
    .B(\u_deb0.Output ),
    .Y(_0561_));
 sg13g2_nor3_1 _2353_ (.A(net172),
    .B(net440),
    .C(_0561_),
    .Y(_0114_));
 sg13g2_nor2_2 _2354_ (.A(_0959_),
    .B(net440),
    .Y(_0562_));
 sg13g2_a21oi_1 _2355_ (.A1(net431),
    .A2(_0562_),
    .Y(_0563_),
    .B1(net169));
 sg13g2_o21ai_1 _2356_ (.B1(_0563_),
    .Y(_0564_),
    .A1(net431),
    .A2(_0562_));
 sg13g2_inv_1 _2357_ (.Y(_0115_),
    .A(_0564_));
 sg13g2_a21oi_1 _2358_ (.A1(net431),
    .A2(_0562_),
    .Y(_0565_),
    .B1(net646));
 sg13g2_and3_1 _2359_ (.X(_0566_),
    .A(net646),
    .B(net431),
    .C(_0562_));
 sg13g2_nor3_1 _2360_ (.A(net173),
    .B(_0565_),
    .C(_0566_),
    .Y(_0116_));
 sg13g2_nor2_1 _2361_ (.A(net856),
    .B(_0566_),
    .Y(_0567_));
 sg13g2_and2_1 _2362_ (.A(net856),
    .B(_0566_),
    .X(_0568_));
 sg13g2_nor3_1 _2363_ (.A(net168),
    .B(_0567_),
    .C(_0568_),
    .Y(_0117_));
 sg13g2_nor2_1 _2364_ (.A(net874),
    .B(_0568_),
    .Y(_0569_));
 sg13g2_and2_1 _2365_ (.A(net874),
    .B(_0568_),
    .X(_0570_));
 sg13g2_nor3_1 _2366_ (.A(net168),
    .B(_0569_),
    .C(_0570_),
    .Y(_0118_));
 sg13g2_nor2_1 _2367_ (.A(net831),
    .B(_0570_),
    .Y(_0571_));
 sg13g2_and2_1 _2368_ (.A(net831),
    .B(_0570_),
    .X(_0572_));
 sg13g2_nor3_1 _2369_ (.A(net168),
    .B(net832),
    .C(_0572_),
    .Y(_0119_));
 sg13g2_nor2_1 _2370_ (.A(net869),
    .B(_0572_),
    .Y(_0573_));
 sg13g2_and2_1 _2371_ (.A(net869),
    .B(_0572_),
    .X(_0574_));
 sg13g2_nor3_1 _2372_ (.A(net168),
    .B(_0573_),
    .C(_0574_),
    .Y(_0120_));
 sg13g2_nor2_1 _2373_ (.A(net873),
    .B(_0574_),
    .Y(_0575_));
 sg13g2_and2_1 _2374_ (.A(net873),
    .B(_0574_),
    .X(_0576_));
 sg13g2_nor3_1 _2375_ (.A(net168),
    .B(_0575_),
    .C(_0576_),
    .Y(_0121_));
 sg13g2_a21oi_1 _2376_ (.A1(net885),
    .A2(_0576_),
    .Y(_0577_),
    .B1(net168));
 sg13g2_o21ai_1 _2377_ (.B1(_0577_),
    .Y(_0578_),
    .A1(net885),
    .A2(_0576_));
 sg13g2_inv_1 _2378_ (.Y(_0122_),
    .A(_0578_));
 sg13g2_nor2_1 _2379_ (.A(change1),
    .B(\u_deb1.Output ),
    .Y(_0579_));
 sg13g2_nor3_1 _2380_ (.A(net172),
    .B(net434),
    .C(_0579_),
    .Y(_0123_));
 sg13g2_nor2_2 _2381_ (.A(_0958_),
    .B(net434),
    .Y(_0580_));
 sg13g2_a21oi_1 _2382_ (.A1(net430),
    .A2(_0580_),
    .Y(_0581_),
    .B1(net162));
 sg13g2_o21ai_1 _2383_ (.B1(_0581_),
    .Y(_0582_),
    .A1(net430),
    .A2(_0580_));
 sg13g2_inv_1 _2384_ (.Y(_0124_),
    .A(_0582_));
 sg13g2_a21oi_1 _2385_ (.A1(net430),
    .A2(_0580_),
    .Y(_0583_),
    .B1(net595));
 sg13g2_and3_1 _2386_ (.X(_0584_),
    .A(net595),
    .B(net430),
    .C(_0580_));
 sg13g2_nor3_1 _2387_ (.A(net162),
    .B(_0583_),
    .C(_0584_),
    .Y(_0125_));
 sg13g2_nor2_1 _2388_ (.A(net857),
    .B(_0584_),
    .Y(_0585_));
 sg13g2_and2_1 _2389_ (.A(net857),
    .B(_0584_),
    .X(_0586_));
 sg13g2_nor3_1 _2390_ (.A(net162),
    .B(_0585_),
    .C(_0586_),
    .Y(_0126_));
 sg13g2_nor2_1 _2391_ (.A(net799),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_and2_1 _2392_ (.A(net155),
    .B(_0586_),
    .X(_0588_));
 sg13g2_nor3_1 _2393_ (.A(net162),
    .B(net800),
    .C(_0588_),
    .Y(_0127_));
 sg13g2_nor2_1 _2394_ (.A(net887),
    .B(_0588_),
    .Y(_0589_));
 sg13g2_and2_1 _2395_ (.A(net887),
    .B(_0588_),
    .X(_0590_));
 sg13g2_nor3_1 _2396_ (.A(net162),
    .B(_0589_),
    .C(_0590_),
    .Y(_0128_));
 sg13g2_nor2_1 _2397_ (.A(net860),
    .B(_0590_),
    .Y(_0591_));
 sg13g2_and2_1 _2398_ (.A(net860),
    .B(_0590_),
    .X(_0592_));
 sg13g2_nor3_1 _2399_ (.A(net162),
    .B(net861),
    .C(_0592_),
    .Y(_0129_));
 sg13g2_nor2_1 _2400_ (.A(net853),
    .B(_0592_),
    .Y(_0593_));
 sg13g2_and2_1 _2401_ (.A(net853),
    .B(_0592_),
    .X(_0594_));
 sg13g2_nor3_1 _2402_ (.A(net162),
    .B(net854),
    .C(_0594_),
    .Y(_0130_));
 sg13g2_a21oi_1 _2403_ (.A1(net878),
    .A2(_0594_),
    .Y(_0595_),
    .B1(net162));
 sg13g2_o21ai_1 _2404_ (.B1(_0595_),
    .Y(_0596_),
    .A1(net878),
    .A2(_0594_));
 sg13g2_inv_1 _2405_ (.Y(_0131_),
    .A(_0596_));
 sg13g2_nor2_1 _2406_ (.A(_0959_),
    .B(net173),
    .Y(_0132_));
 sg13g2_nor2_1 _2407_ (.A(change2),
    .B(\u_deb2.Output ),
    .Y(_0597_));
 sg13g2_nor3_1 _2408_ (.A(net172),
    .B(net436),
    .C(_0597_),
    .Y(_0133_));
 sg13g2_nor2_2 _2409_ (.A(_0957_),
    .B(net436),
    .Y(_0598_));
 sg13g2_a21oi_1 _2410_ (.A1(net429),
    .A2(_0598_),
    .Y(_0599_),
    .B1(net161));
 sg13g2_o21ai_1 _2411_ (.B1(_0599_),
    .Y(_0600_),
    .A1(net429),
    .A2(_0598_));
 sg13g2_inv_1 _2412_ (.Y(_0134_),
    .A(_0600_));
 sg13g2_a21oi_1 _2413_ (.A1(net429),
    .A2(_0598_),
    .Y(_0601_),
    .B1(net571));
 sg13g2_and3_1 _2414_ (.X(_0602_),
    .A(net571),
    .B(net429),
    .C(_0598_));
 sg13g2_nor3_1 _2415_ (.A(net161),
    .B(net572),
    .C(_0602_),
    .Y(_0135_));
 sg13g2_nor2_1 _2416_ (.A(net852),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_and2_1 _2417_ (.A(net852),
    .B(_0602_),
    .X(_0604_));
 sg13g2_nor3_1 _2418_ (.A(net161),
    .B(_0603_),
    .C(_0604_),
    .Y(_0136_));
 sg13g2_nor2_1 _2419_ (.A(net880),
    .B(_0604_),
    .Y(_0605_));
 sg13g2_and2_1 _2420_ (.A(net880),
    .B(_0604_),
    .X(_0606_));
 sg13g2_nor3_1 _2421_ (.A(net161),
    .B(_0605_),
    .C(_0606_),
    .Y(_0137_));
 sg13g2_nor2_1 _2422_ (.A(net154),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_and2_1 _2423_ (.A(net154),
    .B(_0606_),
    .X(_0608_));
 sg13g2_nor3_1 _2424_ (.A(net161),
    .B(_0607_),
    .C(_0608_),
    .Y(_0138_));
 sg13g2_nor2_1 _2425_ (.A(net848),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_and2_1 _2426_ (.A(net848),
    .B(_0608_),
    .X(_0610_));
 sg13g2_nor3_1 _2427_ (.A(net161),
    .B(net849),
    .C(_0610_),
    .Y(_0139_));
 sg13g2_nor2_1 _2428_ (.A(net876),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_and2_1 _2429_ (.A(net876),
    .B(_0610_),
    .X(_0612_));
 sg13g2_nor3_1 _2430_ (.A(net161),
    .B(_0611_),
    .C(_0612_),
    .Y(_0140_));
 sg13g2_a21oi_1 _2431_ (.A1(net886),
    .A2(_0612_),
    .Y(_0613_),
    .B1(net161));
 sg13g2_o21ai_1 _2432_ (.B1(_0613_),
    .Y(_0614_),
    .A1(net886),
    .A2(_0612_));
 sg13g2_inv_1 _2433_ (.Y(_0141_),
    .A(_0614_));
 sg13g2_nor2_1 _2434_ (.A(_0958_),
    .B(net172),
    .Y(_0142_));
 sg13g2_nor2_1 _2435_ (.A(change3),
    .B(\u_deb3.Output ),
    .Y(_0615_));
 sg13g2_nor3_1 _2436_ (.A(net172),
    .B(net438),
    .C(_0615_),
    .Y(_0143_));
 sg13g2_nor2_2 _2437_ (.A(_0956_),
    .B(net438),
    .Y(_0616_));
 sg13g2_a21oi_1 _2438_ (.A1(net428),
    .A2(_0616_),
    .Y(_0617_),
    .B1(net169));
 sg13g2_o21ai_1 _2439_ (.B1(_0617_),
    .Y(_0618_),
    .A1(net428),
    .A2(_0616_));
 sg13g2_inv_1 _2440_ (.Y(_0144_),
    .A(_0618_));
 sg13g2_a21oi_1 _2441_ (.A1(net428),
    .A2(_0616_),
    .Y(_0619_),
    .B1(net587));
 sg13g2_and3_1 _2442_ (.X(_0620_),
    .A(net587),
    .B(net428),
    .C(_0616_));
 sg13g2_nor3_1 _2443_ (.A(net169),
    .B(_0619_),
    .C(_0620_),
    .Y(_0145_));
 sg13g2_nor2_1 _2444_ (.A(net875),
    .B(_0620_),
    .Y(_0621_));
 sg13g2_and2_1 _2445_ (.A(net875),
    .B(_0620_),
    .X(_0622_));
 sg13g2_nor3_1 _2446_ (.A(net168),
    .B(_0621_),
    .C(_0622_),
    .Y(_0146_));
 sg13g2_nor2_1 _2447_ (.A(net153),
    .B(_0622_),
    .Y(_0623_));
 sg13g2_and2_1 _2448_ (.A(net153),
    .B(_0622_),
    .X(_0624_));
 sg13g2_nor3_1 _2449_ (.A(net168),
    .B(_0623_),
    .C(_0624_),
    .Y(_0147_));
 sg13g2_nor2_1 _2450_ (.A(net152),
    .B(_0624_),
    .Y(_0625_));
 sg13g2_and2_1 _2451_ (.A(net892),
    .B(_0624_),
    .X(_0626_));
 sg13g2_nor3_1 _2452_ (.A(net169),
    .B(_0625_),
    .C(_0626_),
    .Y(_0148_));
 sg13g2_nor2_1 _2453_ (.A(net870),
    .B(_0626_),
    .Y(_0627_));
 sg13g2_and2_1 _2454_ (.A(net870),
    .B(_0626_),
    .X(_0628_));
 sg13g2_nor3_1 _2455_ (.A(net169),
    .B(net871),
    .C(_0628_),
    .Y(_0149_));
 sg13g2_nor2_1 _2456_ (.A(net151),
    .B(_0628_),
    .Y(_0629_));
 sg13g2_and2_1 _2457_ (.A(net151),
    .B(_0628_),
    .X(_0630_));
 sg13g2_nor3_1 _2458_ (.A(net169),
    .B(_0629_),
    .C(_0630_),
    .Y(_0150_));
 sg13g2_a21oi_1 _2459_ (.A1(net888),
    .A2(_0630_),
    .Y(_0631_),
    .B1(net169));
 sg13g2_o21ai_1 _2460_ (.B1(_0631_),
    .Y(_0632_),
    .A1(net888),
    .A2(_0630_));
 sg13g2_inv_1 _2461_ (.Y(_0151_),
    .A(net889));
 sg13g2_nor2_1 _2462_ (.A(_0957_),
    .B(net172),
    .Y(_0152_));
 sg13g2_nor2_1 _2463_ (.A(_0956_),
    .B(net170),
    .Y(_0153_));
 sg13g2_nor2_1 _2464_ (.A(\u_edge.Output ),
    .B(\u_deb4.Output ),
    .Y(_0633_));
 sg13g2_nor3_1 _2465_ (.A(net170),
    .B(net432),
    .C(_0633_),
    .Y(_0154_));
 sg13g2_or2_1 _2466_ (.X(_0173_),
    .B(net442),
    .A(net452));
 sg13g2_nor4_1 _2467_ (.A(net473),
    .B(net491),
    .C(net453),
    .D(net461),
    .Y(_0634_));
 sg13g2_nand2b_1 _2468_ (.Y(_0159_),
    .B(_0634_),
    .A_N(_0173_));
 sg13g2_nor2_1 _2469_ (.A(_0955_),
    .B(net170),
    .Y(_0160_));
 sg13g2_or2_1 _2470_ (.X(_0163_),
    .B(net465),
    .A(net460));
 sg13g2_or2_1 _2471_ (.X(_0166_),
    .B(net451),
    .A(net467));
 sg13g2_or2_1 _2472_ (.X(_0169_),
    .B(net443),
    .A(net466));
 sg13g2_nor2_1 _2473_ (.A(\u_edge.Output ),
    .B(net590),
    .Y(_0635_));
 sg13g2_nor2_1 _2474_ (.A(net165),
    .B(net591),
    .Y(_0170_));
 sg13g2_nor4_1 _2475_ (.A(net462),
    .B(net472),
    .C(net468),
    .D(net459),
    .Y(_0636_));
 sg13g2_nand2b_1 _2476_ (.Y(_0178_),
    .B(_0636_),
    .A_N(_0163_));
 sg13g2_nor4_1 _2477_ (.A(net444),
    .B(net496),
    .C(net448),
    .D(net454),
    .Y(_0637_));
 sg13g2_nand2b_1 _2478_ (.Y(_0183_),
    .B(_0637_),
    .A_N(_0166_));
 sg13g2_nor4_1 _2479_ (.A(net458),
    .B(net471),
    .C(net455),
    .D(net447),
    .Y(_0638_));
 sg13g2_nand2b_1 _2480_ (.Y(_0188_),
    .B(_0638_),
    .A_N(_0169_));
 sg13g2_nand2b_2 _2481_ (.Y(_0639_),
    .B(net149),
    .A_N(net148));
 sg13g2_nor2_2 _2482_ (.A(_1063_),
    .B(_0639_),
    .Y(_0640_));
 sg13g2_and2_1 _2483_ (.A(_1077_),
    .B(_0640_),
    .X(_0641_));
 sg13g2_nand2_2 _2484_ (.Y(_0642_),
    .A(net836),
    .B(net895));
 sg13g2_nand3_1 _2485_ (.B(net836),
    .C(net895),
    .A(net149),
    .Y(_0643_));
 sg13g2_nor2_1 _2486_ (.A(net148),
    .B(_0643_),
    .Y(_0644_));
 sg13g2_and2_1 _2487_ (.A(_1077_),
    .B(_0644_),
    .X(_0645_));
 sg13g2_a22oi_1 _2488_ (.Y(_0646_),
    .B1(_0645_),
    .B2(\ascii3[0] ),
    .A2(_0641_),
    .A1(\ascii3[16] ));
 sg13g2_nor4_2 _2489_ (.A(\u_uart.rom.addr[7] ),
    .B(\u_uart.rom.addr[6] ),
    .C(\u_uart.rom.addr[5] ),
    .Y(_0647_),
    .D(\u_uart.rom.addr[4] ));
 sg13g2_and2_1 _2490_ (.A(_1076_),
    .B(_0647_),
    .X(_0648_));
 sg13g2_nand2_1 _2491_ (.Y(_0649_),
    .A(_1076_),
    .B(_0647_));
 sg13g2_nor2_1 _2492_ (.A(net147),
    .B(net149),
    .Y(_0650_));
 sg13g2_or2_1 _2493_ (.X(_0651_),
    .B(\u_uart.rom.addr[0] ),
    .A(\u_uart.rom.addr[1] ));
 sg13g2_nor3_1 _2494_ (.A(net147),
    .B(net149),
    .C(_0651_),
    .Y(_0652_));
 sg13g2_nor4_2 _2495_ (.A(\u_uart.rom.addr[7] ),
    .B(\u_uart.rom.addr[6] ),
    .C(\u_uart.rom.addr[5] ),
    .Y(_0653_),
    .D(_0937_));
 sg13g2_and2_1 _2496_ (.A(_1076_),
    .B(_0653_),
    .X(_0654_));
 sg13g2_nand2_2 _2497_ (.Y(_0655_),
    .A(_1076_),
    .B(_0653_));
 sg13g2_nand2_2 _2498_ (.Y(_0656_),
    .A(net147),
    .B(net149));
 sg13g2_and4_1 _2499_ (.A(net147),
    .B(net150),
    .C(\u_uart.rom.addr[1] ),
    .D(\u_uart.rom.addr[0] ),
    .X(_0657_));
 sg13g2_a22oi_1 _2500_ (.Y(_0658_),
    .B1(_0654_),
    .B2(_0657_),
    .A2(_0652_),
    .A1(_0648_));
 sg13g2_nor3_1 _2501_ (.A(_1064_),
    .B(_0642_),
    .C(_0649_),
    .Y(_0659_));
 sg13g2_nor2_1 _2502_ (.A(_1079_),
    .B(_0659_),
    .Y(_0660_));
 sg13g2_nor3_1 _2503_ (.A(net149),
    .B(_1063_),
    .C(_0649_),
    .Y(_0661_));
 sg13g2_and2_1 _2504_ (.A(net147),
    .B(_0661_),
    .X(_0662_));
 sg13g2_nor3_2 _2505_ (.A(_1063_),
    .B(_0655_),
    .C(_0656_),
    .Y(_0663_));
 sg13g2_and2_1 _2506_ (.A(\ascii2[0] ),
    .B(_0663_),
    .X(_0664_));
 sg13g2_nand2b_2 _2507_ (.Y(_0665_),
    .B(_0650_),
    .A_N(_0642_));
 sg13g2_nor2_2 _2508_ (.A(_0655_),
    .B(_0665_),
    .Y(_0666_));
 sg13g2_a221oi_1 _2509_ (.B2(\ascii1[0] ),
    .C1(_0664_),
    .B1(_0666_),
    .A1(\ascii0[0] ),
    .Y(_0667_),
    .A2(_0662_));
 sg13g2_nand4_1 _2510_ (.B(_0658_),
    .C(_0660_),
    .A(_0646_),
    .Y(_0668_),
    .D(_0667_));
 sg13g2_o21ai_1 _2511_ (.B1(_0665_),
    .Y(_0669_),
    .A1(_1063_),
    .A2(_0656_));
 sg13g2_nand2b_1 _2512_ (.Y(_0670_),
    .B(_0650_),
    .A_N(_1063_));
 sg13g2_a22oi_1 _2513_ (.Y(_0671_),
    .B1(_0669_),
    .B2(_0647_),
    .A2(_0653_),
    .A1(_0644_));
 sg13g2_o21ai_1 _2514_ (.B1(_0671_),
    .Y(_0672_),
    .A1(_1067_),
    .A2(_0670_));
 sg13g2_a21o_1 _2515_ (.A2(_0672_),
    .A1(_1076_),
    .B1(_0984_),
    .X(_0673_));
 sg13g2_nor2_2 _2516_ (.A(_0655_),
    .B(_0670_),
    .Y(_0674_));
 sg13g2_nand2_1 _2517_ (.Y(_0675_),
    .A(\ascii1[16] ),
    .B(_0674_));
 sg13g2_and2_1 _2518_ (.A(_0644_),
    .B(_0648_),
    .X(_0676_));
 sg13g2_nor3_2 _2519_ (.A(_0651_),
    .B(_0655_),
    .C(_0656_),
    .Y(_0677_));
 sg13g2_a22oi_1 _2520_ (.Y(_0678_),
    .B1(_0677_),
    .B2(\ascii2[8] ),
    .A2(_0676_),
    .A1(\ascii0[16] ));
 sg13g2_nor2_1 _2521_ (.A(_1064_),
    .B(_0651_),
    .Y(_0679_));
 sg13g2_and2_1 _2522_ (.A(_0648_),
    .B(_0679_),
    .X(_0680_));
 sg13g2_nand2_2 _2523_ (.Y(_0681_),
    .A(\u_uart.rom.addr[1] ),
    .B(_0938_));
 sg13g2_nor3_1 _2524_ (.A(net147),
    .B(net149),
    .C(_0681_),
    .Y(_0682_));
 sg13g2_inv_1 _2525_ (.Y(_0683_),
    .A(_0682_));
 sg13g2_nor2_2 _2526_ (.A(_0655_),
    .B(_0683_),
    .Y(_0684_));
 sg13g2_a22oi_1 _2527_ (.Y(_0685_),
    .B1(_0684_),
    .B2(\ascii1[8] ),
    .A2(_0680_),
    .A1(\ascii0[8] ));
 sg13g2_nor3_2 _2528_ (.A(_1064_),
    .B(_0642_),
    .C(_0655_),
    .Y(_0686_));
 sg13g2_nor3_2 _2529_ (.A(_1078_),
    .B(_0639_),
    .C(_0681_),
    .Y(_0687_));
 sg13g2_a22oi_1 _2530_ (.Y(_0688_),
    .B1(_0687_),
    .B2(\ascii3[8] ),
    .A2(_0686_),
    .A1(\ascii2[16] ));
 sg13g2_nand4_1 _2531_ (.B(_0678_),
    .C(_0685_),
    .A(_0675_),
    .Y(_0689_),
    .D(_0688_));
 sg13g2_nor3_1 _2532_ (.A(_0668_),
    .B(_0673_),
    .C(_0689_),
    .Y(_0690_));
 sg13g2_o21ai_1 _2533_ (.B1(net157),
    .Y(_0691_),
    .A1(net776),
    .A2(net146));
 sg13g2_nor2_1 _2534_ (.A(_0690_),
    .B(net777),
    .Y(_0189_));
 sg13g2_nor3_1 _2535_ (.A(_0639_),
    .B(_0655_),
    .C(_0681_),
    .Y(_0692_));
 sg13g2_o21ai_1 _2536_ (.B1(_0683_),
    .Y(_0693_),
    .A1(_0651_),
    .A2(_0656_));
 sg13g2_a22oi_1 _2537_ (.Y(_0694_),
    .B1(_0693_),
    .B2(_0648_),
    .A2(_0652_),
    .A1(_1077_));
 sg13g2_nand2b_1 _2538_ (.Y(_0695_),
    .B(_0694_),
    .A_N(_0692_));
 sg13g2_nand2_1 _2539_ (.Y(_0696_),
    .A(_0640_),
    .B(_0654_));
 sg13g2_nand2_1 _2540_ (.Y(_0697_),
    .A(_1077_),
    .B(_0679_));
 sg13g2_nand3_1 _2541_ (.B(_0696_),
    .C(_0697_),
    .A(net146),
    .Y(_0698_));
 sg13g2_and2_1 _2542_ (.A(\ascii0[1] ),
    .B(_0662_),
    .X(_0699_));
 sg13g2_nand2_1 _2543_ (.Y(_0700_),
    .A(\ascii1[9] ),
    .B(_0684_));
 sg13g2_a22oi_1 _2544_ (.Y(_0701_),
    .B1(_0687_),
    .B2(\ascii3[9] ),
    .A2(_0677_),
    .A1(\ascii2[9] ));
 sg13g2_a22oi_1 _2545_ (.Y(_0702_),
    .B1(_0676_),
    .B2(\ascii0[17] ),
    .A2(_0663_),
    .A1(\ascii2[1] ));
 sg13g2_a22oi_1 _2546_ (.Y(_0703_),
    .B1(_0686_),
    .B2(\ascii2[17] ),
    .A2(_0680_),
    .A1(\ascii0[9] ));
 sg13g2_a22oi_1 _2547_ (.Y(_0704_),
    .B1(_0645_),
    .B2(\ascii3[1] ),
    .A2(_0641_),
    .A1(\ascii3[17] ));
 sg13g2_a22oi_1 _2548_ (.Y(_0705_),
    .B1(_0674_),
    .B2(\ascii1[17] ),
    .A2(_0666_),
    .A1(\ascii1[1] ));
 sg13g2_and4_1 _2549_ (.A(_0702_),
    .B(_0703_),
    .C(_0704_),
    .D(_0705_),
    .X(_0706_));
 sg13g2_nand3_1 _2550_ (.B(_0701_),
    .C(_0706_),
    .A(_0700_),
    .Y(_0707_));
 sg13g2_nor4_1 _2551_ (.A(_0695_),
    .B(_0698_),
    .C(_0699_),
    .D(_0707_),
    .Y(_0708_));
 sg13g2_o21ai_1 _2552_ (.B1(net157),
    .Y(_0709_),
    .A1(net750),
    .A2(net146));
 sg13g2_nor2_1 _2553_ (.A(_0708_),
    .B(net751),
    .Y(_0190_));
 sg13g2_a22oi_1 _2554_ (.Y(_0710_),
    .B1(_0680_),
    .B2(\ascii0[10] ),
    .A2(_0645_),
    .A1(\ascii3[2] ));
 sg13g2_nand2_1 _2555_ (.Y(_0711_),
    .A(\ascii3[10] ),
    .B(_0687_));
 sg13g2_nand3_1 _2556_ (.B(_0710_),
    .C(_0711_),
    .A(_0660_),
    .Y(_0712_));
 sg13g2_a21oi_1 _2557_ (.A1(\ascii0[2] ),
    .A2(_0662_),
    .Y(_0713_),
    .B1(_0712_));
 sg13g2_or2_1 _2558_ (.X(_0714_),
    .B(_0657_),
    .A(_0640_));
 sg13g2_a22oi_1 _2559_ (.Y(_0715_),
    .B1(_0714_),
    .B2(_0648_),
    .A2(_0654_),
    .A1(_1065_));
 sg13g2_o21ai_1 _2560_ (.B1(_0715_),
    .Y(_0716_),
    .A1(_1078_),
    .A2(_0665_));
 sg13g2_nor2_1 _2561_ (.A(_0984_),
    .B(_0716_),
    .Y(_0717_));
 sg13g2_a22oi_1 _2562_ (.Y(_0718_),
    .B1(_0677_),
    .B2(\ascii2[10] ),
    .A2(_0666_),
    .A1(\ascii1[2] ));
 sg13g2_a22oi_1 _2563_ (.Y(_0719_),
    .B1(_0684_),
    .B2(\ascii1[10] ),
    .A2(_0663_),
    .A1(\ascii2[2] ));
 sg13g2_and3_1 _2564_ (.X(_0720_),
    .A(_0717_),
    .B(_0718_),
    .C(_0719_));
 sg13g2_o21ai_1 _2565_ (.B1(net157),
    .Y(_0721_),
    .A1(net795),
    .A2(net146));
 sg13g2_a21oi_1 _2566_ (.A1(_0713_),
    .A2(_0720_),
    .Y(_0191_),
    .B1(_0721_));
 sg13g2_nand2_1 _2567_ (.Y(_0722_),
    .A(_0654_),
    .B(_0679_));
 sg13g2_or2_1 _2568_ (.X(_0723_),
    .B(_0651_),
    .A(_0639_));
 sg13g2_o21ai_1 _2569_ (.B1(_0723_),
    .Y(_0724_),
    .A1(_0656_),
    .A2(_0681_));
 sg13g2_a22oi_1 _2570_ (.Y(_0725_),
    .B1(_0724_),
    .B2(_0648_),
    .A2(_0682_),
    .A1(_1077_));
 sg13g2_nand2_1 _2571_ (.Y(_0726_),
    .A(_0722_),
    .B(_0725_));
 sg13g2_nand3_1 _2572_ (.B(_1080_),
    .C(_0697_),
    .A(net146),
    .Y(_0727_));
 sg13g2_and2_1 _2573_ (.A(\ascii0[3] ),
    .B(_0662_),
    .X(_0728_));
 sg13g2_nand2_1 _2574_ (.Y(_0729_),
    .A(\ascii0[11] ),
    .B(_0680_));
 sg13g2_a22oi_1 _2575_ (.Y(_0730_),
    .B1(_0687_),
    .B2(\ascii3[11] ),
    .A2(_0645_),
    .A1(\ascii3[3] ));
 sg13g2_a22oi_1 _2576_ (.Y(_0731_),
    .B1(_0677_),
    .B2(\ascii2[11] ),
    .A2(_0663_),
    .A1(\ascii2[3] ));
 sg13g2_a22oi_1 _2577_ (.Y(_0732_),
    .B1(_0684_),
    .B2(\ascii1[11] ),
    .A2(_0666_),
    .A1(\ascii1[3] ));
 sg13g2_nand4_1 _2578_ (.B(_0730_),
    .C(_0731_),
    .A(_0729_),
    .Y(_0733_),
    .D(_0732_));
 sg13g2_nor4_1 _2579_ (.A(_0726_),
    .B(_0727_),
    .C(_0728_),
    .D(_0733_),
    .Y(_0734_));
 sg13g2_o21ai_1 _2580_ (.B1(net157),
    .Y(_0735_),
    .A1(net790),
    .A2(net146));
 sg13g2_nor2_1 _2581_ (.A(_0734_),
    .B(net791),
    .Y(_0192_));
 sg13g2_nor3_1 _2582_ (.A(_0645_),
    .B(_0659_),
    .C(_0661_),
    .Y(_0736_));
 sg13g2_o21ai_1 _2583_ (.B1(_0654_),
    .Y(_0737_),
    .A1(_0640_),
    .A2(_0669_));
 sg13g2_nand2_1 _2584_ (.Y(_0738_),
    .A(_0658_),
    .B(_0737_));
 sg13g2_nor4_1 _2585_ (.A(_0645_),
    .B(_0659_),
    .C(_0661_),
    .D(_0738_),
    .Y(_0739_));
 sg13g2_a22oi_1 _2586_ (.Y(_0740_),
    .B1(_0687_),
    .B2(\ascii3[12] ),
    .A2(_0686_),
    .A1(\ascii2[20] ));
 sg13g2_a22oi_1 _2587_ (.Y(_0741_),
    .B1(_0680_),
    .B2(\ascii0[12] ),
    .A2(_0676_),
    .A1(\ascii0[20] ));
 sg13g2_a22oi_1 _2588_ (.Y(_0742_),
    .B1(_0677_),
    .B2(\ascii2[12] ),
    .A2(_0641_),
    .A1(\ascii3[20] ));
 sg13g2_nand3_1 _2589_ (.B(_0741_),
    .C(_0742_),
    .A(_0740_),
    .Y(_0743_));
 sg13g2_a221oi_1 _2590_ (.B2(\ascii1[12] ),
    .C1(_0743_),
    .B1(_0684_),
    .A1(\ascii1[20] ),
    .Y(_0744_),
    .A2(_0674_));
 sg13g2_nand3_1 _2591_ (.B(_0739_),
    .C(_0744_),
    .A(_0717_),
    .Y(_0745_));
 sg13g2_o21ai_1 _2592_ (.B1(_0745_),
    .Y(_0746_),
    .A1(net793),
    .A2(net146));
 sg13g2_nor2_1 _2593_ (.A(net164),
    .B(net794),
    .Y(_0193_));
 sg13g2_nand2_1 _2594_ (.Y(_0747_),
    .A(_1064_),
    .B(_0639_));
 sg13g2_a22oi_1 _2595_ (.Y(_0748_),
    .B1(_0747_),
    .B2(_0647_),
    .A2(_0653_),
    .A1(net147));
 sg13g2_nor3_1 _2596_ (.A(\u_uart.rom.addr[1] ),
    .B(_1067_),
    .C(_0639_),
    .Y(_0749_));
 sg13g2_nor2_1 _2597_ (.A(net148),
    .B(_0651_),
    .Y(_0750_));
 sg13g2_a21oi_1 _2598_ (.A1(_0653_),
    .A2(_0750_),
    .Y(_0751_),
    .B1(_0749_));
 sg13g2_o21ai_1 _2599_ (.B1(_0751_),
    .Y(_0752_),
    .A1(_0681_),
    .A2(_0748_));
 sg13g2_nand2_1 _2600_ (.Y(_0753_),
    .A(_1076_),
    .B(_0752_));
 sg13g2_a21oi_1 _2601_ (.A1(_1076_),
    .A2(_0672_),
    .Y(_0754_),
    .B1(_0687_));
 sg13g2_nand3_1 _2602_ (.B(_0753_),
    .C(_0754_),
    .A(_0736_),
    .Y(_0755_));
 sg13g2_nor2_1 _2603_ (.A(_0677_),
    .B(_0684_),
    .Y(_0756_));
 sg13g2_nor4_1 _2604_ (.A(_0674_),
    .B(_0676_),
    .C(_0680_),
    .D(_0686_),
    .Y(_0757_));
 sg13g2_nand2_1 _2605_ (.Y(_0758_),
    .A(_0756_),
    .B(_0757_));
 sg13g2_nor3_1 _2606_ (.A(_0738_),
    .B(_0755_),
    .C(_0758_),
    .Y(_0759_));
 sg13g2_nor3_1 _2607_ (.A(_0695_),
    .B(_0716_),
    .C(_0726_),
    .Y(_0760_));
 sg13g2_a21oi_1 _2608_ (.A1(_0759_),
    .A2(_0760_),
    .Y(_0761_),
    .B1(_0727_));
 sg13g2_a21oi_1 _2609_ (.A1(net566),
    .A2(_0984_),
    .Y(_0762_),
    .B1(_0761_));
 sg13g2_nor2_1 _2610_ (.A(net164),
    .B(net567),
    .Y(_0194_));
 sg13g2_nor2b_1 _2611_ (.A(_0673_),
    .B_N(_0760_),
    .Y(_0763_));
 sg13g2_o21ai_1 _2612_ (.B1(net157),
    .Y(_0764_),
    .A1(net766),
    .A2(_0983_));
 sg13g2_nor2_1 _2613_ (.A(_0763_),
    .B(net767),
    .Y(_0195_));
 sg13g2_nor2_2 _2614_ (.A(net825),
    .B(net163),
    .Y(_0765_));
 sg13g2_or2_1 _2615_ (.X(_0766_),
    .B(net163),
    .A(\u_uart.uart_tx_inst.state[0] ));
 sg13g2_o21ai_1 _2616_ (.B1(_0977_),
    .Y(_0767_),
    .A1(net561),
    .A2(net541));
 sg13g2_nor3_1 _2617_ (.A(net723),
    .B(net850),
    .C(_0767_),
    .Y(_0768_));
 sg13g2_o21ai_1 _2618_ (.B1(net145),
    .Y(_0769_),
    .A1(net606),
    .A2(_0768_));
 sg13g2_inv_1 _2619_ (.Y(_0196_),
    .A(_0769_));
 sg13g2_nor4_1 _2620_ (.A(change3),
    .B(change2),
    .C(change1),
    .D(net809),
    .Y(_0770_));
 sg13g2_nor2_1 _2621_ (.A(net172),
    .B(net810),
    .Y(_0197_));
 sg13g2_nor3_1 _2622_ (.A(\u_uart.uart_tx_inst.state[2] ),
    .B(net906),
    .C(\u_uart.uart_tx_inst.state[3] ),
    .Y(_0771_));
 sg13g2_or3_1 _2623_ (.A(\u_uart.uart_tx_inst.state[2] ),
    .B(net561),
    .C(\u_uart.uart_tx_inst.state[3] ),
    .X(_0772_));
 sg13g2_and2_1 _2624_ (.A(_0976_),
    .B(_0772_),
    .X(_0773_));
 sg13g2_nor2_1 _2625_ (.A(net759),
    .B(_0773_),
    .Y(_0774_));
 sg13g2_and2_1 _2626_ (.A(net759),
    .B(_0772_),
    .X(_0775_));
 sg13g2_nor3_1 _2627_ (.A(_0766_),
    .B(_0774_),
    .C(_0775_),
    .Y(_0198_));
 sg13g2_nand2b_1 _2628_ (.Y(_0776_),
    .B(_0772_),
    .A_N(_0976_));
 sg13g2_nand2_2 _2629_ (.Y(_0777_),
    .A(net145),
    .B(_0776_));
 sg13g2_nor2_1 _2630_ (.A(net717),
    .B(_0775_),
    .Y(_0778_));
 sg13g2_nand2_2 _2631_ (.Y(_0779_),
    .A(net717),
    .B(net759));
 sg13g2_nor2_2 _2632_ (.A(net140),
    .B(_0779_),
    .Y(_0780_));
 sg13g2_nor3_1 _2633_ (.A(_0777_),
    .B(net718),
    .C(_0780_),
    .Y(_0199_));
 sg13g2_xnor2_1 _2634_ (.Y(_0781_),
    .A(net804),
    .B(_0780_));
 sg13g2_nor2_1 _2635_ (.A(_0777_),
    .B(_0781_),
    .Y(_0200_));
 sg13g2_nand3_1 _2636_ (.B(net804),
    .C(_0780_),
    .A(net883),
    .Y(_0782_));
 sg13g2_a21oi_1 _2637_ (.A1(net804),
    .A2(_0780_),
    .Y(_0783_),
    .B1(net883));
 sg13g2_nor2_1 _2638_ (.A(_0777_),
    .B(_0783_),
    .Y(_0784_));
 sg13g2_and2_1 _2639_ (.A(_0782_),
    .B(_0784_),
    .X(_0201_));
 sg13g2_a221oi_1 _2640_ (.B2(_0942_),
    .C1(_0777_),
    .B1(_0782_),
    .A1(_0964_),
    .Y(_0202_),
    .A2(_0780_));
 sg13g2_nor2_1 _2641_ (.A(_0963_),
    .B(_0779_),
    .Y(_0785_));
 sg13g2_nor2_1 _2642_ (.A(_0965_),
    .B(_0779_),
    .Y(_0786_));
 sg13g2_inv_1 _2643_ (.Y(_0787_),
    .A(_0786_));
 sg13g2_a22oi_1 _2644_ (.Y(_0788_),
    .B1(_0773_),
    .B2(_0787_),
    .A2(net140),
    .A1(net780));
 sg13g2_o21ai_1 _2645_ (.B1(net144),
    .Y(_0789_),
    .A1(net780),
    .A2(_0785_));
 sg13g2_nor2_1 _2646_ (.A(_0788_),
    .B(_0789_),
    .Y(_0203_));
 sg13g2_nand3_1 _2647_ (.B(_0772_),
    .C(_0786_),
    .A(net890),
    .Y(_0790_));
 sg13g2_a21oi_1 _2648_ (.A1(_0772_),
    .A2(_0786_),
    .Y(_0791_),
    .B1(net890));
 sg13g2_nor2_1 _2649_ (.A(_0777_),
    .B(_0791_),
    .Y(_0792_));
 sg13g2_and2_1 _2650_ (.A(_0790_),
    .B(_0792_),
    .X(_0204_));
 sg13g2_and3_2 _2651_ (.X(_0793_),
    .A(net842),
    .B(\u_uart.uart_tx_inst.clk_count[6] ),
    .C(_0786_));
 sg13g2_xor2_1 _2652_ (.B(_0790_),
    .A(net842),
    .X(_0794_));
 sg13g2_nor2_1 _2653_ (.A(_0777_),
    .B(net843),
    .Y(_0205_));
 sg13g2_nand2_1 _2654_ (.Y(_0795_),
    .A(net865),
    .B(_0793_));
 sg13g2_a22oi_1 _2655_ (.Y(_0796_),
    .B1(_0773_),
    .B2(_0795_),
    .A2(net140),
    .A1(net865));
 sg13g2_o21ai_1 _2656_ (.B1(net144),
    .Y(_0797_),
    .A1(net865),
    .A2(_0793_));
 sg13g2_nor2_1 _2657_ (.A(net866),
    .B(_0797_),
    .Y(_0206_));
 sg13g2_nand3_1 _2658_ (.B(\u_uart.uart_tx_inst.clk_count[8] ),
    .C(_0793_),
    .A(net640),
    .Y(_0798_));
 sg13g2_a22oi_1 _2659_ (.Y(_0799_),
    .B1(_0773_),
    .B2(_0798_),
    .A2(net140),
    .A1(net640));
 sg13g2_a21oi_1 _2660_ (.A1(\u_uart.uart_tx_inst.clk_count[8] ),
    .A2(_0793_),
    .Y(_0800_),
    .B1(net640));
 sg13g2_nor3_1 _2661_ (.A(_0766_),
    .B(_0799_),
    .C(net641),
    .Y(_0207_));
 sg13g2_nand2b_1 _2662_ (.Y(_0801_),
    .B(_0772_),
    .A_N(_0798_));
 sg13g2_a21oi_1 _2663_ (.A1(_0941_),
    .A2(_0801_),
    .Y(_0208_),
    .B1(_0777_));
 sg13g2_and3_1 _2664_ (.X(_0209_),
    .A(net486),
    .B(net142),
    .C(net138));
 sg13g2_and3_1 _2665_ (.X(_0210_),
    .A(net478),
    .B(net142),
    .C(net138));
 sg13g2_and3_1 _2666_ (.X(_0211_),
    .A(net512),
    .B(net143),
    .C(net139));
 sg13g2_and3_1 _2667_ (.X(_0212_),
    .A(net474),
    .B(net142),
    .C(net138));
 sg13g2_and3_1 _2668_ (.X(_0213_),
    .A(net502),
    .B(net142),
    .C(net138));
 sg13g2_and3_1 _2669_ (.X(_0214_),
    .A(net487),
    .B(net142),
    .C(net138));
 sg13g2_and3_1 _2670_ (.X(_0215_),
    .A(net497),
    .B(net142),
    .C(net138));
 sg13g2_and3_1 _2671_ (.X(_0216_),
    .A(net494),
    .B(net144),
    .C(net139));
 sg13g2_and3_1 _2672_ (.X(_0217_),
    .A(net482),
    .B(net144),
    .C(net139));
 sg13g2_and3_1 _2673_ (.X(_0218_),
    .A(net484),
    .B(net144),
    .C(net139));
 sg13g2_and3_1 _2674_ (.X(_0219_),
    .A(net500),
    .B(net144),
    .C(net139));
 sg13g2_and3_1 _2675_ (.X(_0220_),
    .A(net476),
    .B(net145),
    .C(net141));
 sg13g2_and3_1 _2676_ (.X(_0221_),
    .A(net498),
    .B(net145),
    .C(net141));
 sg13g2_and3_1 _2677_ (.X(_0222_),
    .A(net479),
    .B(net145),
    .C(net141));
 sg13g2_and3_1 _2678_ (.X(_0223_),
    .A(net488),
    .B(net145),
    .C(net141));
 sg13g2_and3_1 _2679_ (.X(_0224_),
    .A(net475),
    .B(net143),
    .C(net140));
 sg13g2_and3_1 _2680_ (.X(_0225_),
    .A(net481),
    .B(net143),
    .C(net140));
 sg13g2_and3_1 _2681_ (.X(_0226_),
    .A(net492),
    .B(net143),
    .C(net140));
 sg13g2_and3_1 _2682_ (.X(_0227_),
    .A(net506),
    .B(net143),
    .C(net138));
 sg13g2_and3_1 _2683_ (.X(_0228_),
    .A(net493),
    .B(net142),
    .C(net139));
 sg13g2_and3_1 _2684_ (.X(_0229_),
    .A(net490),
    .B(net142),
    .C(net138));
 sg13g2_nor3_1 _2685_ (.A(_0961_),
    .B(net850),
    .C(_0976_),
    .Y(_0802_));
 sg13g2_and2_1 _2686_ (.A(net884),
    .B(_0802_),
    .X(_0803_));
 sg13g2_o21ai_1 _2687_ (.B1(net145),
    .Y(_0804_),
    .A1(net884),
    .A2(_0802_));
 sg13g2_nor2_1 _2688_ (.A(_0803_),
    .B(_0804_),
    .Y(_0230_));
 sg13g2_and2_1 _2689_ (.A(net862),
    .B(_0803_),
    .X(_0805_));
 sg13g2_o21ai_1 _2690_ (.B1(net145),
    .Y(_0806_),
    .A1(net862),
    .A2(_0803_));
 sg13g2_nor2_1 _2691_ (.A(_0805_),
    .B(_0806_),
    .Y(_0231_));
 sg13g2_o21ai_1 _2692_ (.B1(_0765_),
    .Y(_0807_),
    .A1(net536),
    .A2(_0805_));
 sg13g2_a21oi_1 _2693_ (.A1(net536),
    .A2(_0805_),
    .Y(_0232_),
    .B1(_0807_));
 sg13g2_nor4_1 _2694_ (.A(\u_uart.uart_tx_inst.state[0] ),
    .B(net723),
    .C(\u_uart.uart_tx_inst.state[3] ),
    .D(_0776_),
    .Y(_0808_));
 sg13g2_nand2b_1 _2695_ (.Y(_0809_),
    .B(net728),
    .A_N(_0808_));
 sg13g2_a21oi_1 _2696_ (.A1(_0984_),
    .A2(net729),
    .Y(_0233_),
    .B1(net163));
 sg13g2_nand2b_1 _2697_ (.Y(_0810_),
    .B(\u_uart.uart_tx_inst.bit_index[0] ),
    .A_N(\u_uart.uart_tx_inst.tx_data[5] ));
 sg13g2_o21ai_1 _2698_ (.B1(_0810_),
    .Y(_0811_),
    .A1(\u_uart.uart_tx_inst.bit_index[0] ),
    .A2(\u_uart.uart_tx_inst.tx_data[4] ));
 sg13g2_nand3b_1 _2699_ (.B(\u_uart.uart_tx_inst.tx_data[6] ),
    .C(\u_uart.uart_tx_inst.bit_index[1] ),
    .Y(_0812_),
    .A_N(\u_uart.uart_tx_inst.bit_index[0] ));
 sg13g2_mux4_1 _2700_ (.S0(\u_uart.uart_tx_inst.bit_index[0] ),
    .A0(\u_uart.uart_tx_inst.tx_data[0] ),
    .A1(\u_uart.uart_tx_inst.tx_data[1] ),
    .A2(\u_uart.uart_tx_inst.tx_data[2] ),
    .A3(\u_uart.uart_tx_inst.tx_data[3] ),
    .S1(\u_uart.uart_tx_inst.bit_index[1] ),
    .X(_0813_));
 sg13g2_nand2b_1 _2701_ (.Y(_0814_),
    .B(_0813_),
    .A_N(net536));
 sg13g2_o21ai_1 _2702_ (.B1(_0812_),
    .Y(_0815_),
    .A1(\u_uart.uart_tx_inst.bit_index[1] ),
    .A2(_0811_));
 sg13g2_a21oi_1 _2703_ (.A1(net536),
    .A2(_0815_),
    .Y(_0816_),
    .B1(_0961_));
 sg13g2_nand2_1 _2704_ (.Y(_0817_),
    .A(_0814_),
    .B(_0816_));
 sg13g2_a21oi_1 _2705_ (.A1(_0940_),
    .A2(net141),
    .Y(_0818_),
    .B1(\u_uart.uart_tx_inst.state[3] ));
 sg13g2_a21oi_1 _2706_ (.A1(_0817_),
    .A2(_0818_),
    .Y(_0819_),
    .B1(net825));
 sg13g2_nor2_1 _2707_ (.A(net163),
    .B(net826),
    .Y(_0234_));
 sg13g2_a221oi_1 _2708_ (.B2(net548),
    .C1(net166),
    .B1(_1082_),
    .A1(_0939_),
    .Y(_0235_),
    .A2(_0987_));
 sg13g2_nor3_1 _2709_ (.A(\u_uart.state[0] ),
    .B(\u_uart.state[3] ),
    .C(\u_uart.state[1] ),
    .Y(_0820_));
 sg13g2_or2_1 _2710_ (.X(_0821_),
    .B(_0820_),
    .A(_0962_));
 sg13g2_a21oi_1 _2711_ (.A1(\u_uart.state[1] ),
    .A2(_1079_),
    .Y(_0822_),
    .B1(_0821_));
 sg13g2_nand2_2 _2712_ (.Y(_0823_),
    .A(_0986_),
    .B(_0822_));
 sg13g2_nor2_1 _2713_ (.A(_1081_),
    .B(_0821_),
    .Y(_0824_));
 sg13g2_or2_1 _2714_ (.X(_0825_),
    .B(_0821_),
    .A(_1081_));
 sg13g2_o21ai_1 _2715_ (.B1(net157),
    .Y(_0826_),
    .A1(_0938_),
    .A2(net125));
 sg13g2_a21oi_1 _2716_ (.A1(_0938_),
    .A2(net118),
    .Y(_0236_),
    .B1(_0826_));
 sg13g2_nand2_1 _2717_ (.Y(_0827_),
    .A(net836),
    .B(net125));
 sg13g2_nand3_1 _2718_ (.B(_0651_),
    .C(net119),
    .A(_0642_),
    .Y(_0828_));
 sg13g2_a21oi_1 _2719_ (.A1(_0827_),
    .A2(_0828_),
    .Y(_0237_),
    .B1(net166));
 sg13g2_xnor2_1 _2720_ (.Y(_0829_),
    .A(net150),
    .B(_0642_));
 sg13g2_a22oi_1 _2721_ (.Y(_0830_),
    .B1(net119),
    .B2(_0829_),
    .A2(net125),
    .A1(net150));
 sg13g2_nor2_1 _2722_ (.A(net171),
    .B(_0830_),
    .Y(_0238_));
 sg13g2_xnor2_1 _2723_ (.Y(_0831_),
    .A(net148),
    .B(_0643_));
 sg13g2_a22oi_1 _2724_ (.Y(_0832_),
    .B1(net119),
    .B2(_0831_),
    .A2(net125),
    .A1(net148));
 sg13g2_nor2_1 _2725_ (.A(net171),
    .B(_0832_),
    .Y(_0239_));
 sg13g2_and2_1 _2726_ (.A(net864),
    .B(_0657_),
    .X(_0833_));
 sg13g2_xnor2_1 _2727_ (.Y(_0834_),
    .A(_0937_),
    .B(_0657_));
 sg13g2_a22oi_1 _2728_ (.Y(_0835_),
    .B1(net119),
    .B2(_0834_),
    .A2(net127),
    .A1(net864));
 sg13g2_nor2_1 _2729_ (.A(net171),
    .B(_0835_),
    .Y(_0240_));
 sg13g2_xor2_1 _2730_ (.B(_0833_),
    .A(net891),
    .X(_0836_));
 sg13g2_a22oi_1 _2731_ (.Y(_0837_),
    .B1(net121),
    .B2(_0836_),
    .A2(net127),
    .A1(net891));
 sg13g2_nor2_1 _2732_ (.A(net171),
    .B(_0837_),
    .Y(_0241_));
 sg13g2_nand4_1 _2733_ (.B(net905),
    .C(net864),
    .A(net756),
    .Y(_0838_),
    .D(_0657_));
 sg13g2_a22oi_1 _2734_ (.Y(_0839_),
    .B1(net119),
    .B2(_0838_),
    .A2(net125),
    .A1(net756));
 sg13g2_a21oi_1 _2735_ (.A1(\u_uart.rom.addr[5] ),
    .A2(_0833_),
    .Y(_0840_),
    .B1(net756));
 sg13g2_nor3_1 _2736_ (.A(net171),
    .B(_0839_),
    .C(net757),
    .Y(_0242_));
 sg13g2_nand2_1 _2737_ (.Y(_0841_),
    .A(net815),
    .B(net125));
 sg13g2_nor2_2 _2738_ (.A(_0936_),
    .B(_0838_),
    .Y(_0842_));
 sg13g2_nand2b_1 _2739_ (.Y(_0843_),
    .B(net119),
    .A_N(_0842_));
 sg13g2_a221oi_1 _2740_ (.B2(_0843_),
    .C1(net171),
    .B1(_0841_),
    .A1(_0936_),
    .Y(_0243_),
    .A2(_0838_));
 sg13g2_nand2_1 _2741_ (.Y(_0844_),
    .A(net877),
    .B(_0842_));
 sg13g2_a22oi_1 _2742_ (.Y(_0845_),
    .B1(net119),
    .B2(_0844_),
    .A2(net125),
    .A1(net877));
 sg13g2_o21ai_1 _2743_ (.B1(net159),
    .Y(_0846_),
    .A1(net877),
    .A2(_0842_));
 sg13g2_nor2_1 _2744_ (.A(_0845_),
    .B(_0846_),
    .Y(_0244_));
 sg13g2_nor4_1 _2745_ (.A(_0934_),
    .B(_0935_),
    .C(_0936_),
    .D(_0838_),
    .Y(_0847_));
 sg13g2_nand3_1 _2746_ (.B(\u_uart.rom.addr[8] ),
    .C(_0842_),
    .A(net637),
    .Y(_0848_));
 sg13g2_a22oi_1 _2747_ (.Y(_0849_),
    .B1(net119),
    .B2(_0848_),
    .A2(net125),
    .A1(net637));
 sg13g2_a21oi_1 _2748_ (.A1(\u_uart.rom.addr[8] ),
    .A2(_0842_),
    .Y(_0850_),
    .B1(net637));
 sg13g2_nor3_1 _2749_ (.A(net171),
    .B(_0849_),
    .C(net638),
    .Y(_0245_));
 sg13g2_and2_1 _2750_ (.A(net748),
    .B(_0847_),
    .X(_0851_));
 sg13g2_inv_1 _2751_ (.Y(_0852_),
    .A(_0851_));
 sg13g2_a22oi_1 _2752_ (.Y(_0853_),
    .B1(net121),
    .B2(_0852_),
    .A2(net127),
    .A1(net748));
 sg13g2_nor2_1 _2753_ (.A(net748),
    .B(_0847_),
    .Y(_0854_));
 sg13g2_nor3_1 _2754_ (.A(net170),
    .B(_0853_),
    .C(net749),
    .Y(_0246_));
 sg13g2_nand2_1 _2755_ (.Y(_0855_),
    .A(net868),
    .B(_0851_));
 sg13g2_a22oi_1 _2756_ (.Y(_0856_),
    .B1(net120),
    .B2(_0855_),
    .A2(net126),
    .A1(net868));
 sg13g2_o21ai_1 _2757_ (.B1(net158),
    .Y(_0857_),
    .A1(net868),
    .A2(_0851_));
 sg13g2_nor2_1 _2758_ (.A(_0856_),
    .B(_0857_),
    .Y(_0247_));
 sg13g2_nand4_1 _2759_ (.B(net868),
    .C(net748),
    .A(net613),
    .Y(_0858_),
    .D(_0847_));
 sg13g2_a22oi_1 _2760_ (.Y(_0859_),
    .B1(net120),
    .B2(_0858_),
    .A2(net126),
    .A1(net613));
 sg13g2_a21oi_1 _2761_ (.A1(\u_uart.rom.addr[11] ),
    .A2(_0851_),
    .Y(_0860_),
    .B1(net613));
 sg13g2_nor3_1 _2762_ (.A(net170),
    .B(_0859_),
    .C(net614),
    .Y(_0248_));
 sg13g2_nand2_1 _2763_ (.Y(_0861_),
    .A(net611),
    .B(net126));
 sg13g2_nor2_2 _2764_ (.A(_0933_),
    .B(_0858_),
    .Y(_0862_));
 sg13g2_nand2b_1 _2765_ (.Y(_0863_),
    .B(net120),
    .A_N(_0862_));
 sg13g2_a221oi_1 _2766_ (.B2(_0863_),
    .C1(net170),
    .B1(_0861_),
    .A1(_0933_),
    .Y(_0249_),
    .A2(_0858_));
 sg13g2_nand2_1 _2767_ (.Y(_0864_),
    .A(net881),
    .B(_0862_));
 sg13g2_a22oi_1 _2768_ (.Y(_0865_),
    .B1(net120),
    .B2(_0864_),
    .A2(net127),
    .A1(net881));
 sg13g2_o21ai_1 _2769_ (.B1(net160),
    .Y(_0866_),
    .A1(net881),
    .A2(_0862_));
 sg13g2_nor2_1 _2770_ (.A(_0865_),
    .B(_0866_),
    .Y(_0250_));
 sg13g2_nor4_1 _2771_ (.A(_0931_),
    .B(_0932_),
    .C(_0933_),
    .D(_0858_),
    .Y(_0867_));
 sg13g2_nand3_1 _2772_ (.B(\u_uart.rom.addr[14] ),
    .C(_0862_),
    .A(net597),
    .Y(_0868_));
 sg13g2_a22oi_1 _2773_ (.Y(_0869_),
    .B1(net120),
    .B2(_0868_),
    .A2(net126),
    .A1(net597));
 sg13g2_a21oi_1 _2774_ (.A1(\u_uart.rom.addr[14] ),
    .A2(_0862_),
    .Y(_0870_),
    .B1(net597));
 sg13g2_nor3_1 _2775_ (.A(net170),
    .B(_0869_),
    .C(net598),
    .Y(_0251_));
 sg13g2_nand2_1 _2776_ (.Y(_0871_),
    .A(net687),
    .B(net126));
 sg13g2_nor2_2 _2777_ (.A(_0930_),
    .B(_0868_),
    .Y(_0872_));
 sg13g2_nand2b_1 _2778_ (.Y(_0873_),
    .B(net120),
    .A_N(_0872_));
 sg13g2_a221oi_1 _2779_ (.B2(_0873_),
    .C1(net170),
    .B1(_0871_),
    .A1(_0930_),
    .Y(_0252_),
    .A2(_0868_));
 sg13g2_nand2_1 _2780_ (.Y(_0874_),
    .A(net858),
    .B(_0872_));
 sg13g2_a22oi_1 _2781_ (.Y(_0875_),
    .B1(net120),
    .B2(_0874_),
    .A2(net126),
    .A1(net858));
 sg13g2_o21ai_1 _2782_ (.B1(net158),
    .Y(_0876_),
    .A1(net858),
    .A2(_0872_));
 sg13g2_nor2_1 _2783_ (.A(_0875_),
    .B(_0876_),
    .Y(_0253_));
 sg13g2_nand4_1 _2784_ (.B(\u_uart.rom.addr[17] ),
    .C(net687),
    .A(net592),
    .Y(_0877_),
    .D(_0867_));
 sg13g2_a22oi_1 _2785_ (.Y(_0878_),
    .B1(net120),
    .B2(_0877_),
    .A2(net126),
    .A1(net592));
 sg13g2_a21oi_1 _2786_ (.A1(\u_uart.rom.addr[17] ),
    .A2(_0872_),
    .Y(_0879_),
    .B1(net592));
 sg13g2_nor3_1 _2787_ (.A(net165),
    .B(_0878_),
    .C(net593),
    .Y(_0254_));
 sg13g2_or2_1 _2788_ (.X(_0880_),
    .B(_0877_),
    .A(_0929_));
 sg13g2_a22oi_1 _2789_ (.Y(_0881_),
    .B1(net122),
    .B2(_0880_),
    .A2(net126),
    .A1(net774));
 sg13g2_a21oi_1 _2790_ (.A1(_0929_),
    .A2(_0877_),
    .Y(_0882_),
    .B1(net165));
 sg13g2_nor2b_1 _2791_ (.A(_0881_),
    .B_N(_0882_),
    .Y(_0255_));
 sg13g2_nand2_1 _2792_ (.Y(_0883_),
    .A(_0928_),
    .B(_0880_));
 sg13g2_nor2_1 _2793_ (.A(_0928_),
    .B(_0880_),
    .Y(_0884_));
 sg13g2_nor2_1 _2794_ (.A(_0825_),
    .B(_0884_),
    .Y(_0885_));
 sg13g2_a22oi_1 _2795_ (.Y(_0886_),
    .B1(_0883_),
    .B2(_0885_),
    .A2(net124),
    .A1(net761));
 sg13g2_nor2_1 _2796_ (.A(net165),
    .B(_0886_),
    .Y(_0256_));
 sg13g2_nor4_2 _2797_ (.A(_0927_),
    .B(_0928_),
    .C(_0929_),
    .Y(_0887_),
    .D(_0877_));
 sg13g2_o21ai_1 _2798_ (.B1(net122),
    .Y(_0888_),
    .A1(net744),
    .A2(_0884_));
 sg13g2_nor2_1 _2799_ (.A(_0887_),
    .B(_0888_),
    .Y(_0889_));
 sg13g2_a21oi_1 _2800_ (.A1(net744),
    .A2(net124),
    .Y(_0890_),
    .B1(_0889_));
 sg13g2_nor2_1 _2801_ (.A(net166),
    .B(net745),
    .Y(_0257_));
 sg13g2_and2_1 _2802_ (.A(net779),
    .B(_0887_),
    .X(_0891_));
 sg13g2_o21ai_1 _2803_ (.B1(net122),
    .Y(_0892_),
    .A1(net779),
    .A2(_0887_));
 sg13g2_nor2_1 _2804_ (.A(_0891_),
    .B(_0892_),
    .Y(_0893_));
 sg13g2_a21oi_1 _2805_ (.A1(net779),
    .A2(net124),
    .Y(_0894_),
    .B1(_0893_));
 sg13g2_nor2_1 _2806_ (.A(net165),
    .B(_0894_),
    .Y(_0258_));
 sg13g2_nand2_1 _2807_ (.Y(_0895_),
    .A(net735),
    .B(net123));
 sg13g2_a21oi_1 _2808_ (.A1(net735),
    .A2(_0891_),
    .Y(_0896_),
    .B1(_0825_));
 sg13g2_o21ai_1 _2809_ (.B1(_0896_),
    .Y(_0897_),
    .A1(net735),
    .A2(_0891_));
 sg13g2_a21oi_1 _2810_ (.A1(_0895_),
    .A2(_0897_),
    .Y(_0259_),
    .B1(net165));
 sg13g2_a21oi_1 _2811_ (.A1(net735),
    .A2(_0891_),
    .Y(_0898_),
    .B1(net820));
 sg13g2_nand4_1 _2812_ (.B(net735),
    .C(net779),
    .A(net820),
    .Y(_0899_),
    .D(_0887_));
 sg13g2_nor2_1 _2813_ (.A(net118),
    .B(_0898_),
    .Y(_0900_));
 sg13g2_a22oi_1 _2814_ (.Y(_0901_),
    .B1(_0899_),
    .B2(_0900_),
    .A2(net123),
    .A1(net820));
 sg13g2_nor2_1 _2815_ (.A(net165),
    .B(_0901_),
    .Y(_0260_));
 sg13g2_nand2_1 _2816_ (.Y(_0902_),
    .A(_0926_),
    .B(_0899_));
 sg13g2_nor2_2 _2817_ (.A(_0926_),
    .B(_0899_),
    .Y(_0903_));
 sg13g2_nor2_1 _2818_ (.A(net118),
    .B(_0903_),
    .Y(_0904_));
 sg13g2_a22oi_1 _2819_ (.Y(_0905_),
    .B1(_0902_),
    .B2(_0904_),
    .A2(net123),
    .A1(net762));
 sg13g2_nor2_1 _2820_ (.A(net164),
    .B(net763),
    .Y(_0261_));
 sg13g2_nand2_1 _2821_ (.Y(_0906_),
    .A(net786),
    .B(net123));
 sg13g2_a21oi_1 _2822_ (.A1(net786),
    .A2(_0903_),
    .Y(_0907_),
    .B1(net118));
 sg13g2_o21ai_1 _2823_ (.B1(_0907_),
    .Y(_0908_),
    .A1(net786),
    .A2(_0903_));
 sg13g2_a21oi_1 _2824_ (.A1(_0906_),
    .A2(_0908_),
    .Y(_0262_),
    .B1(net164));
 sg13g2_a21oi_1 _2825_ (.A1(net786),
    .A2(_0903_),
    .Y(_0909_),
    .B1(net824));
 sg13g2_nand3_1 _2826_ (.B(net786),
    .C(_0903_),
    .A(net824),
    .Y(_0910_));
 sg13g2_nor2_1 _2827_ (.A(net118),
    .B(_0909_),
    .Y(_0911_));
 sg13g2_a22oi_1 _2828_ (.Y(_0912_),
    .B1(_0910_),
    .B2(_0911_),
    .A2(net123),
    .A1(net824));
 sg13g2_nor2_1 _2829_ (.A(net164),
    .B(_0912_),
    .Y(_0263_));
 sg13g2_nand2b_1 _2830_ (.Y(_0913_),
    .B(_0910_),
    .A_N(net772));
 sg13g2_and4_1 _2831_ (.A(net772),
    .B(\u_uart.rom.addr[27] ),
    .C(\u_uart.rom.addr[26] ),
    .D(_0903_),
    .X(_0914_));
 sg13g2_nor2_1 _2832_ (.A(net118),
    .B(_0914_),
    .Y(_0915_));
 sg13g2_a22oi_1 _2833_ (.Y(_0916_),
    .B1(_0913_),
    .B2(_0915_),
    .A2(net123),
    .A1(net772));
 sg13g2_nor2_1 _2834_ (.A(net164),
    .B(net773),
    .Y(_0264_));
 sg13g2_a21oi_1 _2835_ (.A1(net782),
    .A2(_0914_),
    .Y(_0917_),
    .B1(net118));
 sg13g2_a21oi_1 _2836_ (.A1(net782),
    .A2(net123),
    .Y(_0918_),
    .B1(_0917_));
 sg13g2_o21ai_1 _2837_ (.B1(net158),
    .Y(_0919_),
    .A1(net782),
    .A2(_0914_));
 sg13g2_nor2_1 _2838_ (.A(_0918_),
    .B(_0919_),
    .Y(_0265_));
 sg13g2_and3_1 _2839_ (.X(_0920_),
    .A(net782),
    .B(net122),
    .C(_0914_));
 sg13g2_nor2_1 _2840_ (.A(net769),
    .B(_0920_),
    .Y(_0921_));
 sg13g2_nor2_1 _2841_ (.A(net769),
    .B(net118),
    .Y(_0922_));
 sg13g2_nor3_1 _2842_ (.A(net123),
    .B(_0917_),
    .C(_0922_),
    .Y(_0923_));
 sg13g2_nor3_1 _2843_ (.A(net165),
    .B(net770),
    .C(_0923_),
    .Y(_0266_));
 sg13g2_a21oi_1 _2844_ (.A1(net769),
    .A2(_0920_),
    .Y(_0924_),
    .B1(net879));
 sg13g2_a21oi_1 _2845_ (.A1(net879),
    .A2(_0923_),
    .Y(_0925_),
    .B1(_0924_));
 sg13g2_and2_1 _2846_ (.A(net158),
    .B(_0925_),
    .X(_0267_));
 sg13g2_buf_1 _2847_ (.A(net491),
    .X(_0155_));
 sg13g2_buf_1 _2848_ (.A(net473),
    .X(_0156_));
 sg13g2_buf_1 _2849_ (.A(net461),
    .X(_0157_));
 sg13g2_buf_1 _2850_ (.A(net453),
    .X(_0158_));
 sg13g2_buf_1 _2851_ (.A(net465),
    .X(_0161_));
 sg13g2_buf_1 _2852_ (.A(net460),
    .X(_0162_));
 sg13g2_buf_1 _2853_ (.A(net451),
    .X(_0164_));
 sg13g2_buf_1 _2854_ (.A(net467),
    .X(_0165_));
 sg13g2_buf_1 _2855_ (.A(net443),
    .X(_0167_));
 sg13g2_buf_1 _2856_ (.A(net466),
    .X(_0168_));
 sg13g2_buf_1 _2857_ (.A(net442),
    .X(_0171_));
 sg13g2_buf_1 _2858_ (.A(net452),
    .X(_0172_));
 sg13g2_buf_1 _2859_ (.A(net472),
    .X(_0174_));
 sg13g2_buf_1 _2860_ (.A(net462),
    .X(_0175_));
 sg13g2_buf_1 _2861_ (.A(net459),
    .X(_0176_));
 sg13g2_buf_1 _2862_ (.A(net468),
    .X(_0177_));
 sg13g2_buf_1 _2863_ (.A(net496),
    .X(_0179_));
 sg13g2_buf_1 _2864_ (.A(net444),
    .X(_0180_));
 sg13g2_buf_1 _2865_ (.A(net454),
    .X(_0181_));
 sg13g2_buf_1 _2866_ (.A(net448),
    .X(_0182_));
 sg13g2_buf_1 _2867_ (.A(net471),
    .X(_0184_));
 sg13g2_buf_1 _2868_ (.A(net458),
    .X(_0185_));
 sg13g2_buf_1 _2869_ (.A(net447),
    .X(_0186_));
 sg13g2_buf_1 _2870_ (.A(net455),
    .X(_0187_));
 sg13g2_dfrbpq_2 _2871_ (.RESET_B(net239),
    .D(net446),
    .Q(\u_deb0.counter[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _2872_ (.RESET_B(net105),
    .D(_0010_),
    .Q(\u_deb0.counter[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2873_ (.RESET_B(net103),
    .D(net586),
    .Q(\u_deb0.counter[2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2874_ (.RESET_B(net101),
    .D(net636),
    .Q(\u_deb0.counter[3] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2875_ (.RESET_B(net99),
    .D(_0013_),
    .Q(\u_deb0.counter[4] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _2876_ (.RESET_B(net97),
    .D(net521),
    .Q(\u_deb0.counter[5] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2877_ (.RESET_B(net95),
    .D(net545),
    .Q(\u_deb0.counter[6] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2878_ (.RESET_B(net93),
    .D(_0016_),
    .Q(\u_deb0.counter[7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2879_ (.RESET_B(net91),
    .D(net726),
    .Q(\u_deb0.counter[8] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2880_ (.RESET_B(net89),
    .D(_0018_),
    .Q(\u_deb0.counter[9] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2881_ (.RESET_B(net87),
    .D(net605),
    .Q(\u_deb0.counter[10] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_2 _2882_ (.RESET_B(net85),
    .D(net785),
    .Q(\u_deb0.counter[11] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2883_ (.RESET_B(net83),
    .D(net645),
    .Q(\u_deb0.counter[12] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2884_ (.RESET_B(net81),
    .D(_0022_),
    .Q(\u_deb0.counter[13] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2885_ (.RESET_B(net79),
    .D(_0023_),
    .Q(\u_deb0.counter[14] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2886_ (.RESET_B(net77),
    .D(net823),
    .Q(\u_deb0.counter[15] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2887_ (.RESET_B(net75),
    .D(net678),
    .Q(\u_deb0.counter[16] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2888_ (.RESET_B(net73),
    .D(net553),
    .Q(\u_deb0.counter[17] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2889_ (.RESET_B(net71),
    .D(net511),
    .Q(\u_deb0.counter[18] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2890_ (.RESET_B(net69),
    .D(net31),
    .Q(\u_deb0.counter[19] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _2891_ (.RESET_B(net67),
    .D(net734),
    .Q(\u_deb0.Output ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _2892_ (.RESET_B(net65),
    .D(net464),
    .Q(\u_deb1.counter[0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2893_ (.RESET_B(net63),
    .D(net713),
    .Q(\u_deb1.counter[1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2894_ (.RESET_B(net61),
    .D(net582),
    .Q(\u_deb1.counter[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2895_ (.RESET_B(net59),
    .D(net621),
    .Q(\u_deb1.counter[3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2896_ (.RESET_B(net57),
    .D(net711),
    .Q(\u_deb1.counter[4] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _2897_ (.RESET_B(net55),
    .D(net514),
    .Q(\u_deb1.counter[5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2898_ (.RESET_B(net53),
    .D(net540),
    .Q(\u_deb1.counter[6] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2899_ (.RESET_B(net51),
    .D(net618),
    .Q(\u_deb1.counter[7] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2900_ (.RESET_B(net49),
    .D(net694),
    .Q(\u_deb1.counter[8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2901_ (.RESET_B(net47),
    .D(net698),
    .Q(\u_deb1.counter[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2902_ (.RESET_B(net45),
    .D(net684),
    .Q(\u_deb1.counter[10] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _2903_ (.RESET_B(net43),
    .D(net789),
    .Q(\u_deb1.counter[11] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2904_ (.RESET_B(net41),
    .D(net630),
    .Q(\u_deb1.counter[12] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2905_ (.RESET_B(net39),
    .D(_0043_),
    .Q(\u_deb1.counter[13] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2906_ (.RESET_B(net37),
    .D(net808),
    .Q(\u_deb1.counter[14] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2907_ (.RESET_B(net35),
    .D(_0045_),
    .Q(\u_deb1.counter[15] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2908_ (.RESET_B(net33),
    .D(net755),
    .Q(\u_deb1.counter[16] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2909_ (.RESET_B(net406),
    .D(net547),
    .Q(\u_deb1.counter[17] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2910_ (.RESET_B(net404),
    .D(net526),
    .Q(\u_deb1.counter[18] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2911_ (.RESET_B(net402),
    .D(net30),
    .Q(\u_deb1.counter[19] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2912_ (.RESET_B(net400),
    .D(_0050_),
    .Q(\u_deb1.Output ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _2913_ (.RESET_B(net398),
    .D(net470),
    .Q(\u_deb2.counter[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _2914_ (.RESET_B(net396),
    .D(_0052_),
    .Q(\u_deb2.counter[1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2915_ (.RESET_B(net394),
    .D(net576),
    .Q(\u_deb2.counter[2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2916_ (.RESET_B(net392),
    .D(net655),
    .Q(\u_deb2.counter[3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2917_ (.RESET_B(net390),
    .D(_0055_),
    .Q(\u_deb2.counter[4] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _2918_ (.RESET_B(net388),
    .D(net516),
    .Q(\u_deb2.counter[5] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2919_ (.RESET_B(net386),
    .D(net560),
    .Q(\u_deb2.counter[6] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2920_ (.RESET_B(net384),
    .D(net652),
    .Q(\u_deb2.counter[7] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2921_ (.RESET_B(net382),
    .D(net691),
    .Q(\u_deb2.counter[8] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2922_ (.RESET_B(net380),
    .D(_0060_),
    .Q(\u_deb2.counter[9] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2923_ (.RESET_B(net378),
    .D(net660),
    .Q(\u_deb2.counter[10] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _2924_ (.RESET_B(net376),
    .D(_0062_),
    .Q(\u_deb2.counter[11] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2925_ (.RESET_B(net374),
    .D(net602),
    .Q(\u_deb2.counter[12] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2926_ (.RESET_B(net372),
    .D(_0064_),
    .Q(\u_deb2.counter[13] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2927_ (.RESET_B(net370),
    .D(_0065_),
    .Q(\u_deb2.counter[14] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2928_ (.RESET_B(net368),
    .D(_0066_),
    .Q(\u_deb2.counter[15] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2929_ (.RESET_B(net366),
    .D(net739),
    .Q(\u_deb2.counter[16] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2930_ (.RESET_B(net364),
    .D(net557),
    .Q(\u_deb2.counter[17] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2931_ (.RESET_B(net362),
    .D(net529),
    .Q(\u_deb2.counter[18] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _2932_ (.RESET_B(net360),
    .D(net29),
    .Q(\u_deb2.counter[19] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2933_ (.RESET_B(net358),
    .D(_0071_),
    .Q(\u_deb2.Output ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2934_ (.RESET_B(net356),
    .D(net457),
    .Q(\u_deb3.counter[0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _2935_ (.RESET_B(net354),
    .D(_0073_),
    .Q(\u_deb3.counter[1] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2936_ (.RESET_B(net352),
    .D(net570),
    .Q(\u_deb3.counter[2] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2937_ (.RESET_B(net350),
    .D(net624),
    .Q(\u_deb3.counter[3] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2938_ (.RESET_B(net348),
    .D(_0076_),
    .Q(\u_deb3.counter[4] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _2939_ (.RESET_B(net346),
    .D(net523),
    .Q(\u_deb3.counter[5] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2940_ (.RESET_B(net344),
    .D(net532),
    .Q(\u_deb3.counter[6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2941_ (.RESET_B(net342),
    .D(net681),
    .Q(\u_deb3.counter[7] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2942_ (.RESET_B(net340),
    .D(_0080_),
    .Q(\u_deb3.counter[8] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2943_ (.RESET_B(net338),
    .D(net666),
    .Q(\u_deb3.counter[9] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2944_ (.RESET_B(net336),
    .D(net708),
    .Q(\u_deb3.counter[10] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _2945_ (.RESET_B(net334),
    .D(_0083_),
    .Q(\u_deb3.counter[11] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2946_ (.RESET_B(net332),
    .D(net610),
    .Q(\u_deb3.counter[12] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2947_ (.RESET_B(net330),
    .D(_0085_),
    .Q(\u_deb3.counter[13] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2948_ (.RESET_B(net328),
    .D(net813),
    .Q(\u_deb3.counter[14] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2949_ (.RESET_B(net322),
    .D(_0087_),
    .Q(\u_deb3.counter[15] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2950_ (.RESET_B(net320),
    .D(net701),
    .Q(\u_deb3.counter[16] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2951_ (.RESET_B(net314),
    .D(net551),
    .Q(\u_deb3.counter[17] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2952_ (.RESET_B(net312),
    .D(net519),
    .Q(\u_deb3.counter[18] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2953_ (.RESET_B(net310),
    .D(net28),
    .Q(\u_deb3.counter[19] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _2954_ (.RESET_B(net304),
    .D(net722),
    .Q(\u_deb3.Output ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _2955_ (.RESET_B(net302),
    .D(net450),
    .Q(\u_deb4.counter[0] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _2956_ (.RESET_B(net296),
    .D(net686),
    .Q(\u_deb4.counter[1] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2957_ (.RESET_B(net294),
    .D(net579),
    .Q(\u_deb4.counter[2] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2958_ (.RESET_B(net292),
    .D(net633),
    .Q(\u_deb4.counter[3] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2959_ (.RESET_B(net290),
    .D(net675),
    .Q(\u_deb4.counter[4] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _2960_ (.RESET_B(net278),
    .D(net508),
    .Q(\u_deb4.counter[5] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2961_ (.RESET_B(net266),
    .D(net535),
    .Q(\u_deb4.counter[6] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2962_ (.RESET_B(net264),
    .D(net663),
    .Q(\u_deb4.counter[7] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2963_ (.RESET_B(net238),
    .D(net672),
    .Q(\u_deb4.counter[8] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2964_ (.RESET_B(net236),
    .D(net669),
    .Q(\u_deb4.counter[9] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2965_ (.RESET_B(net234),
    .D(net627),
    .Q(\u_deb4.counter[10] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _2966_ (.RESET_B(net232),
    .D(_0104_),
    .Q(\u_deb4.counter[11] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2967_ (.RESET_B(net230),
    .D(net649),
    .Q(\u_deb4.counter[12] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2968_ (.RESET_B(net228),
    .D(_0106_),
    .Q(\u_deb4.counter[13] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2969_ (.RESET_B(net226),
    .D(net829),
    .Q(\u_deb4.counter[14] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2970_ (.RESET_B(net224),
    .D(_0108_),
    .Q(\u_deb4.counter[15] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2971_ (.RESET_B(net222),
    .D(net705),
    .Q(\u_deb4.counter[16] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2972_ (.RESET_B(net220),
    .D(net555),
    .Q(\u_deb4.counter[17] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2973_ (.RESET_B(net218),
    .D(net505),
    .Q(\u_deb4.counter[18] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2974_ (.RESET_B(net216),
    .D(net27),
    .Q(\u_deb4.counter[19] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2975_ (.RESET_B(net214),
    .D(_0113_),
    .Q(\u_deb4.Output ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2976_ (.RESET_B(net212),
    .D(net441),
    .Q(change0),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _2977_ (.RESET_B(net210),
    .D(_0115_),
    .Q(\u_cnt0.count[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _2978_ (.RESET_B(net208),
    .D(_0116_),
    .Q(\u_cnt0.count[1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _2979_ (.RESET_B(net206),
    .D(_0117_),
    .Q(\u_cnt0.count[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _2980_ (.RESET_B(net204),
    .D(_0118_),
    .Q(\u_cnt0.count[3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _2981_ (.RESET_B(net202),
    .D(net833),
    .Q(\u_cnt0.count[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _2982_ (.RESET_B(net200),
    .D(_0120_),
    .Q(\u_cnt0.count[5] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _2983_ (.RESET_B(net198),
    .D(_0121_),
    .Q(\u_cnt0.count[6] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _2984_ (.RESET_B(net196),
    .D(_0122_),
    .Q(\u_cnt0.count[7] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2985_ (.RESET_B(net194),
    .D(net435),
    .Q(change1),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _2986_ (.RESET_B(net192),
    .D(_0124_),
    .Q(\u_cnt1.count[0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _2987_ (.RESET_B(net190),
    .D(_0125_),
    .Q(\u_cnt1.count[1] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _2988_ (.RESET_B(net188),
    .D(_0126_),
    .Q(\u_cnt1.count[2] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _2989_ (.RESET_B(net186),
    .D(net801),
    .Q(\u_cnt1.count[3] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _2990_ (.RESET_B(net184),
    .D(_0128_),
    .Q(\u_cnt1.count[4] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _2991_ (.RESET_B(net182),
    .D(_0129_),
    .Q(\u_cnt1.count[5] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _2992_ (.RESET_B(net180),
    .D(net855),
    .Q(\u_cnt1.count[6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _2993_ (.RESET_B(net178),
    .D(_0131_),
    .Q(\u_cnt1.count[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2994_ (.RESET_B(net176),
    .D(_0132_),
    .Q(\u_cnt0.state ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2995_ (.RESET_B(net175),
    .D(net437),
    .Q(change2),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _2996_ (.RESET_B(net117),
    .D(_0134_),
    .Q(\u_cnt2.count[0] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _2997_ (.RESET_B(net115),
    .D(_0135_),
    .Q(\u_cnt2.count[1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _2998_ (.RESET_B(net113),
    .D(_0136_),
    .Q(\u_cnt2.count[2] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _2999_ (.RESET_B(net111),
    .D(_0137_),
    .Q(\u_cnt2.count[3] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _3000_ (.RESET_B(net109),
    .D(_0138_),
    .Q(\u_cnt2.count[4] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _3001_ (.RESET_B(net107),
    .D(_0139_),
    .Q(\u_cnt2.count[5] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _3002_ (.RESET_B(net104),
    .D(_0140_),
    .Q(\u_cnt2.count[6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _3003_ (.RESET_B(net100),
    .D(_0141_),
    .Q(\u_cnt2.count[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _3004_ (.RESET_B(net96),
    .D(_0142_),
    .Q(\u_cnt1.state ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3005_ (.RESET_B(net94),
    .D(net439),
    .Q(change3),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _3006_ (.RESET_B(net90),
    .D(_0144_),
    .Q(\u_cnt3.count[0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _3007_ (.RESET_B(net86),
    .D(_0145_),
    .Q(\u_cnt3.count[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _3008_ (.RESET_B(net82),
    .D(_0146_),
    .Q(\u_cnt3.count[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3009_ (.RESET_B(net78),
    .D(_0147_),
    .Q(\u_cnt3.count[3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3010_ (.RESET_B(net74),
    .D(net893),
    .Q(\u_cnt3.count[4] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _3011_ (.RESET_B(net70),
    .D(net872),
    .Q(\u_cnt3.count[5] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _3012_ (.RESET_B(net66),
    .D(_0150_),
    .Q(\u_cnt3.count[6] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _3013_ (.RESET_B(net62),
    .D(_0151_),
    .Q(\u_cnt3.count[7] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _3014_ (.RESET_B(net58),
    .D(_0152_),
    .Q(\u_cnt2.state ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _3015_ (.RESET_B(net56),
    .D(_0153_),
    .Q(\u_cnt3.state ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3016_ (.RESET_B(net54),
    .D(net433),
    .Q(\u_edge.Output ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3017_ (.RESET_B(net50),
    .D(_0155_),
    .Q(\ascii3[8] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3018_ (.RESET_B(net48),
    .D(_0156_),
    .Q(\ascii3[9] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3019_ (.RESET_B(net46),
    .D(_0157_),
    .Q(\ascii3[10] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3020_ (.RESET_B(net44),
    .D(_0158_),
    .Q(\ascii3[11] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3021_ (.RESET_B(net240),
    .D(_0159_),
    .Q(\ascii3[12] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3022_ (.RESET_B(net241),
    .D(_0002_),
    .Q(\u_uart.state[0] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _3023_ (.RESET_B(net242),
    .D(net716),
    .Q(\u_uart.state[1] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3024_ (.RESET_B(net243),
    .D(net847),
    .Q(\u_uart.state[2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3025_ (.RESET_B(net244),
    .D(net607),
    .Q(\u_uart.state[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3026_ (.RESET_B(net245),
    .D(net431),
    .Q(\u_n2a0.ones[0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3027_ (.RESET_B(net246),
    .D(_0274_),
    .Q(\u_n2a0.ones[1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3028_ (.RESET_B(net247),
    .D(_0275_),
    .Q(\u_n2a0.ones[2] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3029_ (.RESET_B(net248),
    .D(_0276_),
    .Q(\u_n2a0.ones[3] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3030_ (.RESET_B(net249),
    .D(_0270_),
    .Q(\u_n2a0.tens[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3031_ (.RESET_B(net250),
    .D(_0271_),
    .Q(\u_n2a0.tens[1] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3032_ (.RESET_B(net251),
    .D(_0272_),
    .Q(\u_n2a0.tens[2] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3033_ (.RESET_B(net252),
    .D(_0273_),
    .Q(\u_n2a0.tens[3] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3034_ (.RESET_B(net254),
    .D(_0268_),
    .Q(\u_n2a0.hundreds[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3035_ (.RESET_B(net42),
    .D(_0269_),
    .Q(\u_n2a0.hundreds[1] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3036_ (.RESET_B(net255),
    .D(_0160_),
    .Q(\u_edge.state ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3037_ (.RESET_B(net256),
    .D(net430),
    .Q(\u_n2a1.ones[0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3038_ (.RESET_B(net257),
    .D(net596),
    .Q(\u_n2a1.ones[1] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3039_ (.RESET_B(net258),
    .D(_0284_),
    .Q(\u_n2a1.ones[2] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3040_ (.RESET_B(net259),
    .D(_0285_),
    .Q(\u_n2a1.ones[3] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3041_ (.RESET_B(net260),
    .D(_0279_),
    .Q(\u_n2a1.tens[0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3042_ (.RESET_B(net261),
    .D(_0280_),
    .Q(\u_n2a1.tens[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3043_ (.RESET_B(net262),
    .D(_0281_),
    .Q(\u_n2a1.tens[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3044_ (.RESET_B(net263),
    .D(_0282_),
    .Q(\u_n2a1.tens[3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3045_ (.RESET_B(net267),
    .D(_0277_),
    .Q(\u_n2a1.hundreds[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3046_ (.RESET_B(net40),
    .D(_0278_),
    .Q(\u_n2a1.hundreds[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3047_ (.RESET_B(net38),
    .D(_0161_),
    .Q(\ascii0[16] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3048_ (.RESET_B(net36),
    .D(_0162_),
    .Q(\ascii0[17] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3049_ (.RESET_B(net268),
    .D(_0163_),
    .Q(\ascii0[20] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3050_ (.RESET_B(net269),
    .D(net429),
    .Q(\u_n2a2.ones[0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _3051_ (.RESET_B(net270),
    .D(_0292_),
    .Q(\u_n2a2.ones[1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _3052_ (.RESET_B(net271),
    .D(_0293_),
    .Q(\u_n2a2.ones[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3053_ (.RESET_B(net272),
    .D(_0294_),
    .Q(\u_n2a2.ones[3] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3054_ (.RESET_B(net273),
    .D(_0288_),
    .Q(\u_n2a2.tens[0] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3055_ (.RESET_B(net274),
    .D(_0289_),
    .Q(\u_n2a2.tens[1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3056_ (.RESET_B(net275),
    .D(_0290_),
    .Q(\u_n2a2.tens[2] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3057_ (.RESET_B(net276),
    .D(_0291_),
    .Q(\u_n2a2.tens[3] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3058_ (.RESET_B(net280),
    .D(_0286_),
    .Q(\u_n2a2.hundreds[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _3059_ (.RESET_B(net34),
    .D(_0287_),
    .Q(\u_n2a2.hundreds[1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3060_ (.RESET_B(net32),
    .D(_0164_),
    .Q(\ascii1[16] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3061_ (.RESET_B(net405),
    .D(_0165_),
    .Q(\ascii1[17] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3062_ (.RESET_B(net281),
    .D(_0166_),
    .Q(\ascii1[20] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3063_ (.RESET_B(net282),
    .D(net428),
    .Q(\u_n2a3.ones[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _3064_ (.RESET_B(net283),
    .D(_0301_),
    .Q(\u_n2a3.ones[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3065_ (.RESET_B(net284),
    .D(_0302_),
    .Q(\u_n2a3.ones[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3066_ (.RESET_B(net285),
    .D(_0303_),
    .Q(\u_n2a3.ones[3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _3067_ (.RESET_B(net286),
    .D(_0297_),
    .Q(\u_n2a3.tens[0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3068_ (.RESET_B(net287),
    .D(_0298_),
    .Q(\u_n2a3.tens[1] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3069_ (.RESET_B(net288),
    .D(_0299_),
    .Q(\u_n2a3.tens[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3070_ (.RESET_B(net289),
    .D(_0300_),
    .Q(\u_n2a3.tens[3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3071_ (.RESET_B(net297),
    .D(_0295_),
    .Q(\u_n2a3.hundreds[0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3072_ (.RESET_B(net403),
    .D(_0296_),
    .Q(\u_n2a3.hundreds[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3073_ (.RESET_B(net401),
    .D(_0167_),
    .Q(\ascii2[16] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3074_ (.RESET_B(net399),
    .D(_0168_),
    .Q(\ascii2[17] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3075_ (.RESET_B(net397),
    .D(_0169_),
    .Q(\ascii2[20] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3076_ (.RESET_B(net395),
    .D(_0170_),
    .Q(start_sending),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _3077_ (.RESET_B(net393),
    .D(_0171_),
    .Q(\ascii3[16] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _3078_ (.RESET_B(net391),
    .D(_0172_),
    .Q(\ascii3[17] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3079_ (.RESET_B(net298),
    .D(_0173_),
    .Q(\ascii3[20] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3080_ (.RESET_B(net299),
    .D(net415),
    .Q(\ascii0[0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3081_ (.RESET_B(net300),
    .D(net419),
    .Q(\ascii0[1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3082_ (.RESET_B(net306),
    .D(net423),
    .Q(\ascii0[2] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _3083_ (.RESET_B(net389),
    .D(net414),
    .Q(\ascii0[3] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _3084_ (.RESET_B(net387),
    .D(_0174_),
    .Q(\ascii0[8] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _3085_ (.RESET_B(net385),
    .D(_0175_),
    .Q(\ascii0[9] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3086_ (.RESET_B(net383),
    .D(_0176_),
    .Q(\ascii0[10] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3087_ (.RESET_B(net381),
    .D(_0177_),
    .Q(\ascii0[11] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3088_ (.RESET_B(net307),
    .D(_0178_),
    .Q(\ascii0[12] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _3089_ (.RESET_B(net308),
    .D(net421),
    .Q(\ascii1[0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _3090_ (.RESET_B(net309),
    .D(net424),
    .Q(\ascii1[1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3091_ (.RESET_B(net315),
    .D(net426),
    .Q(\ascii1[2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3092_ (.RESET_B(net379),
    .D(net425),
    .Q(\ascii1[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3093_ (.RESET_B(net377),
    .D(_0179_),
    .Q(\ascii1[8] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _3094_ (.RESET_B(net375),
    .D(_0180_),
    .Q(\ascii1[9] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3095_ (.RESET_B(net373),
    .D(_0181_),
    .Q(\ascii1[10] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3096_ (.RESET_B(net371),
    .D(_0182_),
    .Q(\ascii1[11] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3097_ (.RESET_B(net316),
    .D(_0183_),
    .Q(\ascii1[12] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3098_ (.RESET_B(net317),
    .D(net413),
    .Q(\ascii2[0] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3099_ (.RESET_B(net318),
    .D(net412),
    .Q(\ascii2[1] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3100_ (.RESET_B(net324),
    .D(net418),
    .Q(\ascii2[2] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3101_ (.RESET_B(net369),
    .D(net417),
    .Q(\ascii2[3] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3102_ (.RESET_B(net367),
    .D(_0184_),
    .Q(\ascii2[8] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3103_ (.RESET_B(net365),
    .D(_0185_),
    .Q(\ascii2[9] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3104_ (.RESET_B(net363),
    .D(_0186_),
    .Q(\ascii2[10] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3105_ (.RESET_B(net361),
    .D(_0187_),
    .Q(\ascii2[11] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _3106_ (.RESET_B(net325),
    .D(_0188_),
    .Q(\ascii2[12] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _3107_ (.RESET_B(net326),
    .D(net427),
    .Q(\ascii3[0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3108_ (.RESET_B(net327),
    .D(net416),
    .Q(\ascii3[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3109_ (.RESET_B(net407),
    .D(net420),
    .Q(\ascii3[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3110_ (.RESET_B(net359),
    .D(net422),
    .Q(\ascii3[3] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _3111_ (.RESET_B(net357),
    .D(net778),
    .Q(\u_uart.uart_tx_inst.tx_data[0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3112_ (.RESET_B(net353),
    .D(net752),
    .Q(\u_uart.uart_tx_inst.tx_data[1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3113_ (.RESET_B(net349),
    .D(net796),
    .Q(\u_uart.uart_tx_inst.tx_data[2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _3114_ (.RESET_B(net345),
    .D(net792),
    .Q(\u_uart.uart_tx_inst.tx_data[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3115_ (.RESET_B(net341),
    .D(_0193_),
    .Q(\u_uart.uart_tx_inst.tx_data[4] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3116_ (.RESET_B(net337),
    .D(_0194_),
    .Q(\u_uart.uart_tx_inst.tx_data[5] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _3117_ (.RESET_B(net333),
    .D(net768),
    .Q(\u_uart.uart_tx_inst.tx_data[6] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _3118_ (.RESET_B(net329),
    .D(_0196_),
    .Q(o_Tx_Done),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3119_ (.RESET_B(net321),
    .D(_0197_),
    .Q(or4_out),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _3120_ (.RESET_B(net319),
    .D(net760),
    .Q(\u_uart.uart_tx_inst.clk_count[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3121_ (.RESET_B(net311),
    .D(net719),
    .Q(\u_uart.uart_tx_inst.clk_count[1] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _3122_ (.RESET_B(net303),
    .D(net805),
    .Q(\u_uart.uart_tx_inst.clk_count[2] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3123_ (.RESET_B(net295),
    .D(_0201_),
    .Q(\u_uart.uart_tx_inst.clk_count[3] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3124_ (.RESET_B(net291),
    .D(net563),
    .Q(\u_uart.uart_tx_inst.clk_count[4] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3125_ (.RESET_B(net277),
    .D(net781),
    .Q(\u_uart.uart_tx_inst.clk_count[5] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3126_ (.RESET_B(net253),
    .D(_0204_),
    .Q(\u_uart.uart_tx_inst.clk_count[6] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3127_ (.RESET_B(net235),
    .D(_0205_),
    .Q(\u_uart.uart_tx_inst.clk_count[7] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _3128_ (.RESET_B(net231),
    .D(net867),
    .Q(\u_uart.uart_tx_inst.clk_count[8] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3129_ (.RESET_B(net227),
    .D(net642),
    .Q(\u_uart.uart_tx_inst.clk_count[9] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3130_ (.RESET_B(net223),
    .D(net565),
    .Q(\u_uart.uart_tx_inst.clk_count[10] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3131_ (.RESET_B(net219),
    .D(_0209_),
    .Q(\u_uart.uart_tx_inst.clk_count[11] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3132_ (.RESET_B(net215),
    .D(_0210_),
    .Q(\u_uart.uart_tx_inst.clk_count[12] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3133_ (.RESET_B(net211),
    .D(_0211_),
    .Q(\u_uart.uart_tx_inst.clk_count[13] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3134_ (.RESET_B(net207),
    .D(_0212_),
    .Q(\u_uart.uart_tx_inst.clk_count[14] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3135_ (.RESET_B(net203),
    .D(_0213_),
    .Q(\u_uart.uart_tx_inst.clk_count[15] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3136_ (.RESET_B(net199),
    .D(_0214_),
    .Q(\u_uart.uart_tx_inst.clk_count[16] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3137_ (.RESET_B(net195),
    .D(_0215_),
    .Q(\u_uart.uart_tx_inst.clk_count[17] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _3138_ (.RESET_B(net191),
    .D(net495),
    .Q(\u_uart.uart_tx_inst.clk_count[18] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3139_ (.RESET_B(net187),
    .D(net483),
    .Q(\u_uart.uart_tx_inst.clk_count[19] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3140_ (.RESET_B(net183),
    .D(net485),
    .Q(\u_uart.uart_tx_inst.clk_count[20] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3141_ (.RESET_B(net179),
    .D(net501),
    .Q(\u_uart.uart_tx_inst.clk_count[21] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3142_ (.RESET_B(net174),
    .D(net477),
    .Q(\u_uart.uart_tx_inst.clk_count[22] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3143_ (.RESET_B(net114),
    .D(net499),
    .Q(\u_uart.uart_tx_inst.clk_count[23] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3144_ (.RESET_B(net110),
    .D(net480),
    .Q(\u_uart.uart_tx_inst.clk_count[24] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3145_ (.RESET_B(net106),
    .D(net489),
    .Q(\u_uart.uart_tx_inst.clk_count[25] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _3146_ (.RESET_B(net98),
    .D(_0224_),
    .Q(\u_uart.uart_tx_inst.clk_count[26] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3147_ (.RESET_B(net88),
    .D(_0225_),
    .Q(\u_uart.uart_tx_inst.clk_count[27] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _3148_ (.RESET_B(net80),
    .D(_0226_),
    .Q(\u_uart.uart_tx_inst.clk_count[28] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3149_ (.RESET_B(net72),
    .D(_0227_),
    .Q(\u_uart.uart_tx_inst.clk_count[29] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _3150_ (.RESET_B(net64),
    .D(_0228_),
    .Q(\u_uart.uart_tx_inst.clk_count[30] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _3151_ (.RESET_B(net52),
    .D(_0229_),
    .Q(\u_uart.uart_tx_inst.clk_count[31] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _3152_ (.RESET_B(net351),
    .D(_0230_),
    .Q(\u_uart.uart_tx_inst.bit_index[0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _3153_ (.RESET_B(net343),
    .D(_0231_),
    .Q(\u_uart.uart_tx_inst.bit_index[1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _3154_ (.RESET_B(net335),
    .D(net537),
    .Q(\u_uart.uart_tx_inst.bit_index[2] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _3155_ (.RESET_B(net323),
    .D(net730),
    .Q(o_Tx_Active),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3156_ (.RESET_B(net305),
    .D(_0234_),
    .Q(o_Tx_Serial),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _3157_ (.RESET_B(net293),
    .D(net549),
    .Q(\u_uart.uart_tx_inst.i_Tx_Start [0]),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _3158_ (.RESET_B(net265),
    .D(_0236_),
    .Q(\u_uart.rom.addr[0] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _3159_ (.RESET_B(net233),
    .D(net837),
    .Q(\u_uart.rom.addr[1] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _3160_ (.RESET_B(net225),
    .D(_0238_),
    .Q(\u_uart.rom.addr[2] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _3161_ (.RESET_B(net217),
    .D(_0239_),
    .Q(\u_uart.rom.addr[3] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _3162_ (.RESET_B(net209),
    .D(_0240_),
    .Q(\u_uart.rom.addr[4] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _3163_ (.RESET_B(net201),
    .D(_0241_),
    .Q(\u_uart.rom.addr[5] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _3164_ (.RESET_B(net193),
    .D(net758),
    .Q(\u_uart.rom.addr[6] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _3165_ (.RESET_B(net185),
    .D(net816),
    .Q(\u_uart.rom.addr[7] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _3166_ (.RESET_B(net177),
    .D(_0244_),
    .Q(\u_uart.rom.addr[8] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _3167_ (.RESET_B(net112),
    .D(net639),
    .Q(\u_uart.rom.addr[9] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _3168_ (.RESET_B(net102),
    .D(_0246_),
    .Q(\u_uart.rom.addr[10] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _3169_ (.RESET_B(net84),
    .D(_0247_),
    .Q(\u_uart.rom.addr[11] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3170_ (.RESET_B(net68),
    .D(net615),
    .Q(\u_uart.rom.addr[12] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3171_ (.RESET_B(net355),
    .D(net612),
    .Q(\u_uart.rom.addr[13] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _3172_ (.RESET_B(net339),
    .D(_0250_),
    .Q(\u_uart.rom.addr[14] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _3173_ (.RESET_B(net313),
    .D(net599),
    .Q(\u_uart.rom.addr[15] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3174_ (.RESET_B(net279),
    .D(net688),
    .Q(\u_uart.rom.addr[16] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _3175_ (.RESET_B(net229),
    .D(net859),
    .Q(\u_uart.rom.addr[17] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _3176_ (.RESET_B(net213),
    .D(net594),
    .Q(\u_uart.rom.addr[18] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _3177_ (.RESET_B(net197),
    .D(net775),
    .Q(\u_uart.rom.addr[19] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3178_ (.RESET_B(net181),
    .D(_0256_),
    .Q(\u_uart.rom.addr[20] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3179_ (.RESET_B(net108),
    .D(_0257_),
    .Q(\u_uart.rom.addr[21] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _3180_ (.RESET_B(net76),
    .D(_0258_),
    .Q(\u_uart.rom.addr[22] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _3181_ (.RESET_B(net347),
    .D(net736),
    .Q(\u_uart.rom.addr[23] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _3182_ (.RESET_B(net301),
    .D(_0260_),
    .Q(\u_uart.rom.addr[24] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _3183_ (.RESET_B(net221),
    .D(_0261_),
    .Q(\u_uart.rom.addr[25] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _3184_ (.RESET_B(net189),
    .D(net787),
    .Q(\u_uart.rom.addr[26] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _3185_ (.RESET_B(net92),
    .D(_0263_),
    .Q(\u_uart.rom.addr[27] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _3186_ (.RESET_B(net331),
    .D(_0264_),
    .Q(\u_uart.rom.addr[28] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _3187_ (.RESET_B(net205),
    .D(net783),
    .Q(\u_uart.rom.addr[29] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _3188_ (.RESET_B(net60),
    .D(net771),
    .Q(\u_uart.rom.addr[30] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _3189_ (.RESET_B(net408),
    .D(_0267_),
    .Q(\u_uart.rom.addr[31] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _3190_ (.RESET_B(net409),
    .D(net542),
    .Q(\u_uart.uart_tx_inst.state[0] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _3191_ (.RESET_B(net410),
    .D(_0001_),
    .Q(\u_uart.uart_tx_inst.state[1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _3192_ (.RESET_B(net411),
    .D(_0006_),
    .Q(\u_uart.uart_tx_inst.state[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _3193_ (.RESET_B(net237),
    .D(_0007_),
    .Q(\u_uart.uart_tx_inst.state[3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _3194_ (.RESET_B(net116),
    .D(_0008_),
    .Q(\u_uart.uart_tx_inst.state[4] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_tiehi _2908__33 (.L_HI(net33));
 sg13g2_tiehi _3059__34 (.L_HI(net34));
 sg13g2_tiehi _2907__35 (.L_HI(net35));
 sg13g2_tiehi _3048__36 (.L_HI(net36));
 sg13g2_tiehi _2906__37 (.L_HI(net37));
 sg13g2_tiehi _3047__38 (.L_HI(net38));
 sg13g2_tiehi _2905__39 (.L_HI(net39));
 sg13g2_tiehi _3046__40 (.L_HI(net40));
 sg13g2_tiehi _2904__41 (.L_HI(net41));
 sg13g2_tiehi _3035__42 (.L_HI(net42));
 sg13g2_tiehi _2903__43 (.L_HI(net43));
 sg13g2_tiehi _3020__44 (.L_HI(net44));
 sg13g2_tiehi _2902__45 (.L_HI(net45));
 sg13g2_tiehi _3019__46 (.L_HI(net46));
 sg13g2_tiehi _2901__47 (.L_HI(net47));
 sg13g2_tiehi _3018__48 (.L_HI(net48));
 sg13g2_tiehi _2900__49 (.L_HI(net49));
 sg13g2_tiehi _3017__50 (.L_HI(net50));
 sg13g2_tiehi _2899__51 (.L_HI(net51));
 sg13g2_tiehi _3151__52 (.L_HI(net52));
 sg13g2_tiehi _2898__53 (.L_HI(net53));
 sg13g2_tiehi _3016__54 (.L_HI(net54));
 sg13g2_tiehi _2897__55 (.L_HI(net55));
 sg13g2_tiehi _3015__56 (.L_HI(net56));
 sg13g2_tiehi _2896__57 (.L_HI(net57));
 sg13g2_tiehi _3014__58 (.L_HI(net58));
 sg13g2_tiehi _2895__59 (.L_HI(net59));
 sg13g2_tiehi _3188__60 (.L_HI(net60));
 sg13g2_tiehi _2894__61 (.L_HI(net61));
 sg13g2_tiehi _3013__62 (.L_HI(net62));
 sg13g2_tiehi _2893__63 (.L_HI(net63));
 sg13g2_tiehi _3150__64 (.L_HI(net64));
 sg13g2_tiehi _2892__65 (.L_HI(net65));
 sg13g2_tiehi _3012__66 (.L_HI(net66));
 sg13g2_tiehi _2891__67 (.L_HI(net67));
 sg13g2_tiehi _3170__68 (.L_HI(net68));
 sg13g2_tiehi _2890__69 (.L_HI(net69));
 sg13g2_tiehi _3011__70 (.L_HI(net70));
 sg13g2_tiehi _2889__71 (.L_HI(net71));
 sg13g2_tiehi _3149__72 (.L_HI(net72));
 sg13g2_tiehi _2888__73 (.L_HI(net73));
 sg13g2_tiehi _3010__74 (.L_HI(net74));
 sg13g2_tiehi _2887__75 (.L_HI(net75));
 sg13g2_tiehi _3180__76 (.L_HI(net76));
 sg13g2_tiehi _2886__77 (.L_HI(net77));
 sg13g2_tiehi _3009__78 (.L_HI(net78));
 sg13g2_tiehi _2885__79 (.L_HI(net79));
 sg13g2_tiehi _3148__80 (.L_HI(net80));
 sg13g2_tiehi _2884__81 (.L_HI(net81));
 sg13g2_tiehi _3008__82 (.L_HI(net82));
 sg13g2_tiehi _2883__83 (.L_HI(net83));
 sg13g2_tiehi _3169__84 (.L_HI(net84));
 sg13g2_tiehi _2882__85 (.L_HI(net85));
 sg13g2_tiehi _3007__86 (.L_HI(net86));
 sg13g2_tiehi _2881__87 (.L_HI(net87));
 sg13g2_tiehi _3147__88 (.L_HI(net88));
 sg13g2_tiehi _2880__89 (.L_HI(net89));
 sg13g2_tiehi _3006__90 (.L_HI(net90));
 sg13g2_tiehi _2879__91 (.L_HI(net91));
 sg13g2_tiehi _3185__92 (.L_HI(net92));
 sg13g2_tiehi _2878__93 (.L_HI(net93));
 sg13g2_tiehi _3005__94 (.L_HI(net94));
 sg13g2_tiehi _2877__95 (.L_HI(net95));
 sg13g2_tiehi _3004__96 (.L_HI(net96));
 sg13g2_tiehi _2876__97 (.L_HI(net97));
 sg13g2_tiehi _3146__98 (.L_HI(net98));
 sg13g2_tiehi _2875__99 (.L_HI(net99));
 sg13g2_tiehi _3003__100 (.L_HI(net100));
 sg13g2_tiehi _2874__101 (.L_HI(net101));
 sg13g2_tiehi _3168__102 (.L_HI(net102));
 sg13g2_tiehi _2873__103 (.L_HI(net103));
 sg13g2_tiehi _3002__104 (.L_HI(net104));
 sg13g2_tiehi _2872__105 (.L_HI(net105));
 sg13g2_tiehi _3145__106 (.L_HI(net106));
 sg13g2_tiehi _3001__107 (.L_HI(net107));
 sg13g2_tiehi _3179__108 (.L_HI(net108));
 sg13g2_tiehi _3000__109 (.L_HI(net109));
 sg13g2_tiehi _3144__110 (.L_HI(net110));
 sg13g2_tiehi _2999__111 (.L_HI(net111));
 sg13g2_tiehi _3167__112 (.L_HI(net112));
 sg13g2_tiehi _2998__113 (.L_HI(net113));
 sg13g2_tiehi _3143__114 (.L_HI(net114));
 sg13g2_tiehi _2997__115 (.L_HI(net115));
 sg13g2_tiehi _3194__116 (.L_HI(net116));
 sg13g2_tiehi _2996__117 (.L_HI(net117));
 sg13g2_tiehi _3142__118 (.L_HI(net174));
 sg13g2_tiehi _2995__119 (.L_HI(net175));
 sg13g2_tiehi _2994__120 (.L_HI(net176));
 sg13g2_tiehi _3166__121 (.L_HI(net177));
 sg13g2_tiehi _2993__122 (.L_HI(net178));
 sg13g2_tiehi _3141__123 (.L_HI(net179));
 sg13g2_tiehi _2992__124 (.L_HI(net180));
 sg13g2_tiehi _3178__125 (.L_HI(net181));
 sg13g2_tiehi _2991__126 (.L_HI(net182));
 sg13g2_tiehi _3140__127 (.L_HI(net183));
 sg13g2_tiehi _2990__128 (.L_HI(net184));
 sg13g2_tiehi _3165__129 (.L_HI(net185));
 sg13g2_tiehi _2989__130 (.L_HI(net186));
 sg13g2_tiehi _3139__131 (.L_HI(net187));
 sg13g2_tiehi _2988__132 (.L_HI(net188));
 sg13g2_tiehi _3184__133 (.L_HI(net189));
 sg13g2_tiehi _2987__134 (.L_HI(net190));
 sg13g2_tiehi _3138__135 (.L_HI(net191));
 sg13g2_tiehi _2986__136 (.L_HI(net192));
 sg13g2_tiehi _3164__137 (.L_HI(net193));
 sg13g2_tiehi _2985__138 (.L_HI(net194));
 sg13g2_tiehi _3137__139 (.L_HI(net195));
 sg13g2_tiehi _2984__140 (.L_HI(net196));
 sg13g2_tiehi _3177__141 (.L_HI(net197));
 sg13g2_tiehi _2983__142 (.L_HI(net198));
 sg13g2_tiehi _3136__143 (.L_HI(net199));
 sg13g2_tiehi _2982__144 (.L_HI(net200));
 sg13g2_tiehi _3163__145 (.L_HI(net201));
 sg13g2_tiehi _2981__146 (.L_HI(net202));
 sg13g2_tiehi _3135__147 (.L_HI(net203));
 sg13g2_tiehi _2980__148 (.L_HI(net204));
 sg13g2_tiehi _3187__149 (.L_HI(net205));
 sg13g2_tiehi _2979__150 (.L_HI(net206));
 sg13g2_tiehi _3134__151 (.L_HI(net207));
 sg13g2_tiehi _2978__152 (.L_HI(net208));
 sg13g2_tiehi _3162__153 (.L_HI(net209));
 sg13g2_tiehi _2977__154 (.L_HI(net210));
 sg13g2_tiehi _3133__155 (.L_HI(net211));
 sg13g2_tiehi _2976__156 (.L_HI(net212));
 sg13g2_tiehi _3176__157 (.L_HI(net213));
 sg13g2_tiehi _2975__158 (.L_HI(net214));
 sg13g2_tiehi _3132__159 (.L_HI(net215));
 sg13g2_tiehi _2974__160 (.L_HI(net216));
 sg13g2_tiehi _3161__161 (.L_HI(net217));
 sg13g2_tiehi _2973__162 (.L_HI(net218));
 sg13g2_tiehi _3131__163 (.L_HI(net219));
 sg13g2_tiehi _2972__164 (.L_HI(net220));
 sg13g2_tiehi _3183__165 (.L_HI(net221));
 sg13g2_tiehi _2971__166 (.L_HI(net222));
 sg13g2_tiehi _3130__167 (.L_HI(net223));
 sg13g2_tiehi _2970__168 (.L_HI(net224));
 sg13g2_tiehi _3160__169 (.L_HI(net225));
 sg13g2_tiehi _2969__170 (.L_HI(net226));
 sg13g2_tiehi _3129__171 (.L_HI(net227));
 sg13g2_tiehi _2968__172 (.L_HI(net228));
 sg13g2_tiehi _3175__173 (.L_HI(net229));
 sg13g2_tiehi _2967__174 (.L_HI(net230));
 sg13g2_tiehi _3128__175 (.L_HI(net231));
 sg13g2_tiehi _2966__176 (.L_HI(net232));
 sg13g2_tiehi _3159__177 (.L_HI(net233));
 sg13g2_tiehi _2965__178 (.L_HI(net234));
 sg13g2_tiehi _3127__179 (.L_HI(net235));
 sg13g2_tiehi _2964__180 (.L_HI(net236));
 sg13g2_tiehi _3193__181 (.L_HI(net237));
 sg13g2_tiehi _2963__182 (.L_HI(net238));
 sg13g2_tiehi _2871__183 (.L_HI(net239));
 sg13g2_tiehi _3021__184 (.L_HI(net240));
 sg13g2_tiehi _3022__185 (.L_HI(net241));
 sg13g2_tiehi _3023__186 (.L_HI(net242));
 sg13g2_tiehi _3024__187 (.L_HI(net243));
 sg13g2_tiehi _3025__188 (.L_HI(net244));
 sg13g2_tiehi _3026__189 (.L_HI(net245));
 sg13g2_tiehi _3027__190 (.L_HI(net246));
 sg13g2_tiehi _3028__191 (.L_HI(net247));
 sg13g2_tiehi _3029__192 (.L_HI(net248));
 sg13g2_tiehi _3030__193 (.L_HI(net249));
 sg13g2_tiehi _3031__194 (.L_HI(net250));
 sg13g2_tiehi _3032__195 (.L_HI(net251));
 sg13g2_tiehi _3033__196 (.L_HI(net252));
 sg13g2_tiehi _3126__197 (.L_HI(net253));
 sg13g2_tiehi _3034__198 (.L_HI(net254));
 sg13g2_tiehi _3036__199 (.L_HI(net255));
 sg13g2_tiehi _3037__200 (.L_HI(net256));
 sg13g2_tiehi _3038__201 (.L_HI(net257));
 sg13g2_tiehi _3039__202 (.L_HI(net258));
 sg13g2_tiehi _3040__203 (.L_HI(net259));
 sg13g2_tiehi _3041__204 (.L_HI(net260));
 sg13g2_tiehi _3042__205 (.L_HI(net261));
 sg13g2_tiehi _3043__206 (.L_HI(net262));
 sg13g2_tiehi _3044__207 (.L_HI(net263));
 sg13g2_tiehi _2962__208 (.L_HI(net264));
 sg13g2_tiehi _3158__209 (.L_HI(net265));
 sg13g2_tiehi _2961__210 (.L_HI(net266));
 sg13g2_tiehi _3045__211 (.L_HI(net267));
 sg13g2_tiehi _3049__212 (.L_HI(net268));
 sg13g2_tiehi _3050__213 (.L_HI(net269));
 sg13g2_tiehi _3051__214 (.L_HI(net270));
 sg13g2_tiehi _3052__215 (.L_HI(net271));
 sg13g2_tiehi _3053__216 (.L_HI(net272));
 sg13g2_tiehi _3054__217 (.L_HI(net273));
 sg13g2_tiehi _3055__218 (.L_HI(net274));
 sg13g2_tiehi _3056__219 (.L_HI(net275));
 sg13g2_tiehi _3057__220 (.L_HI(net276));
 sg13g2_tiehi _3125__221 (.L_HI(net277));
 sg13g2_tiehi _2960__222 (.L_HI(net278));
 sg13g2_tiehi _3174__223 (.L_HI(net279));
 sg13g2_tiehi _3058__224 (.L_HI(net280));
 sg13g2_tiehi _3062__225 (.L_HI(net281));
 sg13g2_tiehi _3063__226 (.L_HI(net282));
 sg13g2_tiehi _3064__227 (.L_HI(net283));
 sg13g2_tiehi _3065__228 (.L_HI(net284));
 sg13g2_tiehi _3066__229 (.L_HI(net285));
 sg13g2_tiehi _3067__230 (.L_HI(net286));
 sg13g2_tiehi _3068__231 (.L_HI(net287));
 sg13g2_tiehi _3069__232 (.L_HI(net288));
 sg13g2_tiehi _3070__233 (.L_HI(net289));
 sg13g2_tiehi _2959__234 (.L_HI(net290));
 sg13g2_tiehi _3124__235 (.L_HI(net291));
 sg13g2_tiehi _2958__236 (.L_HI(net292));
 sg13g2_tiehi _3157__237 (.L_HI(net293));
 sg13g2_tiehi _2957__238 (.L_HI(net294));
 sg13g2_tiehi _3123__239 (.L_HI(net295));
 sg13g2_tiehi _2956__240 (.L_HI(net296));
 sg13g2_tiehi _3071__241 (.L_HI(net297));
 sg13g2_tiehi _3079__242 (.L_HI(net298));
 sg13g2_tiehi _3080__243 (.L_HI(net299));
 sg13g2_tiehi _3081__244 (.L_HI(net300));
 sg13g2_tiehi _3182__245 (.L_HI(net301));
 sg13g2_tiehi _2955__246 (.L_HI(net302));
 sg13g2_tiehi _3122__247 (.L_HI(net303));
 sg13g2_tiehi _2954__248 (.L_HI(net304));
 sg13g2_tiehi _3156__249 (.L_HI(net305));
 sg13g2_tiehi _3082__250 (.L_HI(net306));
 sg13g2_tiehi _3088__251 (.L_HI(net307));
 sg13g2_tiehi _3089__252 (.L_HI(net308));
 sg13g2_tiehi _3090__253 (.L_HI(net309));
 sg13g2_tiehi _2953__254 (.L_HI(net310));
 sg13g2_tiehi _3121__255 (.L_HI(net311));
 sg13g2_tiehi _2952__256 (.L_HI(net312));
 sg13g2_tiehi _3173__257 (.L_HI(net313));
 sg13g2_tiehi _2951__258 (.L_HI(net314));
 sg13g2_tiehi _3091__259 (.L_HI(net315));
 sg13g2_tiehi _3097__260 (.L_HI(net316));
 sg13g2_tiehi _3098__261 (.L_HI(net317));
 sg13g2_tiehi _3099__262 (.L_HI(net318));
 sg13g2_tiehi _3120__263 (.L_HI(net319));
 sg13g2_tiehi _2950__264 (.L_HI(net320));
 sg13g2_tiehi _3119__265 (.L_HI(net321));
 sg13g2_tiehi _2949__266 (.L_HI(net322));
 sg13g2_tiehi _3155__267 (.L_HI(net323));
 sg13g2_tiehi _3100__268 (.L_HI(net324));
 sg13g2_tiehi _3106__269 (.L_HI(net325));
 sg13g2_tiehi _3107__270 (.L_HI(net326));
 sg13g2_tiehi _3108__271 (.L_HI(net327));
 sg13g2_tiehi _2948__272 (.L_HI(net328));
 sg13g2_tiehi _3118__273 (.L_HI(net329));
 sg13g2_tiehi _2947__274 (.L_HI(net330));
 sg13g2_tiehi _3186__275 (.L_HI(net331));
 sg13g2_tiehi _2946__276 (.L_HI(net332));
 sg13g2_tiehi _3117__277 (.L_HI(net333));
 sg13g2_tiehi _2945__278 (.L_HI(net334));
 sg13g2_tiehi _3154__279 (.L_HI(net335));
 sg13g2_tiehi _2944__280 (.L_HI(net336));
 sg13g2_tiehi _3116__281 (.L_HI(net337));
 sg13g2_tiehi _2943__282 (.L_HI(net338));
 sg13g2_tiehi _3172__283 (.L_HI(net339));
 sg13g2_tiehi _2942__284 (.L_HI(net340));
 sg13g2_tiehi _3115__285 (.L_HI(net341));
 sg13g2_tiehi _2941__286 (.L_HI(net342));
 sg13g2_tiehi _3153__287 (.L_HI(net343));
 sg13g2_tiehi _2940__288 (.L_HI(net344));
 sg13g2_tiehi _3114__289 (.L_HI(net345));
 sg13g2_tiehi _2939__290 (.L_HI(net346));
 sg13g2_tiehi _3181__291 (.L_HI(net347));
 sg13g2_tiehi _2938__292 (.L_HI(net348));
 sg13g2_tiehi _3113__293 (.L_HI(net349));
 sg13g2_tiehi _2937__294 (.L_HI(net350));
 sg13g2_tiehi _3152__295 (.L_HI(net351));
 sg13g2_tiehi _2936__296 (.L_HI(net352));
 sg13g2_tiehi _3112__297 (.L_HI(net353));
 sg13g2_tiehi _2935__298 (.L_HI(net354));
 sg13g2_tiehi _3171__299 (.L_HI(net355));
 sg13g2_tiehi _2934__300 (.L_HI(net356));
 sg13g2_tiehi _3111__301 (.L_HI(net357));
 sg13g2_tiehi _2933__302 (.L_HI(net358));
 sg13g2_tiehi _3110__303 (.L_HI(net359));
 sg13g2_tiehi _2932__304 (.L_HI(net360));
 sg13g2_tiehi _3105__305 (.L_HI(net361));
 sg13g2_tiehi _2931__306 (.L_HI(net362));
 sg13g2_tiehi _3104__307 (.L_HI(net363));
 sg13g2_tiehi _2930__308 (.L_HI(net364));
 sg13g2_tiehi _3103__309 (.L_HI(net365));
 sg13g2_tiehi _2929__310 (.L_HI(net366));
 sg13g2_tiehi _3102__311 (.L_HI(net367));
 sg13g2_tiehi _2928__312 (.L_HI(net368));
 sg13g2_tiehi _3101__313 (.L_HI(net369));
 sg13g2_tiehi _2927__314 (.L_HI(net370));
 sg13g2_tiehi _3096__315 (.L_HI(net371));
 sg13g2_tiehi _2926__316 (.L_HI(net372));
 sg13g2_tiehi _3095__317 (.L_HI(net373));
 sg13g2_tiehi _2925__318 (.L_HI(net374));
 sg13g2_tiehi _3094__319 (.L_HI(net375));
 sg13g2_tiehi _2924__320 (.L_HI(net376));
 sg13g2_tiehi _3093__321 (.L_HI(net377));
 sg13g2_tiehi _2923__322 (.L_HI(net378));
 sg13g2_tiehi _3092__323 (.L_HI(net379));
 sg13g2_tiehi _2922__324 (.L_HI(net380));
 sg13g2_tiehi _3087__325 (.L_HI(net381));
 sg13g2_tiehi _2921__326 (.L_HI(net382));
 sg13g2_tiehi _3086__327 (.L_HI(net383));
 sg13g2_tiehi _2920__328 (.L_HI(net384));
 sg13g2_tiehi _3085__329 (.L_HI(net385));
 sg13g2_tiehi _2919__330 (.L_HI(net386));
 sg13g2_tiehi _3084__331 (.L_HI(net387));
 sg13g2_tiehi _2918__332 (.L_HI(net388));
 sg13g2_tiehi _3083__333 (.L_HI(net389));
 sg13g2_tiehi _2917__334 (.L_HI(net390));
 sg13g2_tiehi _3078__335 (.L_HI(net391));
 sg13g2_tiehi _2916__336 (.L_HI(net392));
 sg13g2_tiehi _3077__337 (.L_HI(net393));
 sg13g2_tiehi _2915__338 (.L_HI(net394));
 sg13g2_tiehi _3076__339 (.L_HI(net395));
 sg13g2_tiehi _2914__340 (.L_HI(net396));
 sg13g2_tiehi _3075__341 (.L_HI(net397));
 sg13g2_tiehi _2913__342 (.L_HI(net398));
 sg13g2_tiehi _3074__343 (.L_HI(net399));
 sg13g2_tiehi _2912__344 (.L_HI(net400));
 sg13g2_tiehi _3073__345 (.L_HI(net401));
 sg13g2_tiehi _2911__346 (.L_HI(net402));
 sg13g2_tiehi _3072__347 (.L_HI(net403));
 sg13g2_tiehi _2910__348 (.L_HI(net404));
 sg13g2_tiehi _3061__349 (.L_HI(net405));
 sg13g2_tiehi _2909__350 (.L_HI(net406));
 sg13g2_tiehi _3109__351 (.L_HI(net407));
 sg13g2_tiehi _3189__352 (.L_HI(net408));
 sg13g2_tiehi _3190__353 (.L_HI(net409));
 sg13g2_tiehi _3191__354 (.L_HI(net410));
 sg13g2_tiehi _3192__355 (.L_HI(net411));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_piggy_top_7 (.L_LO(net7));
 sg13g2_tielo tt_um_piggy_top_8 (.L_LO(net8));
 sg13g2_tielo tt_um_piggy_top_9 (.L_LO(net9));
 sg13g2_tielo tt_um_piggy_top_10 (.L_LO(net10));
 sg13g2_tielo tt_um_piggy_top_11 (.L_LO(net11));
 sg13g2_tielo tt_um_piggy_top_12 (.L_LO(net12));
 sg13g2_tielo tt_um_piggy_top_13 (.L_LO(net13));
 sg13g2_tielo tt_um_piggy_top_14 (.L_LO(net14));
 sg13g2_tielo tt_um_piggy_top_15 (.L_LO(net15));
 sg13g2_tielo tt_um_piggy_top_16 (.L_LO(net16));
 sg13g2_tielo tt_um_piggy_top_17 (.L_LO(net17));
 sg13g2_tielo tt_um_piggy_top_18 (.L_LO(net18));
 sg13g2_tielo tt_um_piggy_top_19 (.L_LO(net19));
 sg13g2_tielo tt_um_piggy_top_20 (.L_LO(net20));
 sg13g2_tielo tt_um_piggy_top_21 (.L_LO(net21));
 sg13g2_tielo tt_um_piggy_top_22 (.L_LO(net22));
 sg13g2_tielo tt_um_piggy_top_23 (.L_LO(net23));
 sg13g2_tielo tt_um_piggy_top_24 (.L_LO(net24));
 sg13g2_tielo tt_um_piggy_top_25 (.L_LO(net25));
 sg13g2_tielo tt_um_piggy_top_26 (.L_LO(net26));
 sg13g2_tielo _2974__27 (.L_LO(net27));
 sg13g2_tielo _2953__28 (.L_LO(net28));
 sg13g2_tielo _2932__29 (.L_LO(net29));
 sg13g2_tielo _2911__30 (.L_LO(net30));
 sg13g2_tielo _2890__31 (.L_LO(net31));
 sg13g2_tiehi _3060__32 (.L_HI(net32));
 sg13g2_buf_2 _3545_ (.A(o_Tx_Active),
    .X(uo_out[0]));
 sg13g2_buf_2 _3546_ (.A(o_Tx_Done),
    .X(uo_out[1]));
 sg13g2_buf_8 _3547_ (.A(o_Tx_Serial),
    .X(uo_out[2]));
 sg13g2_buf_8 fanout118 (.A(_0825_),
    .X(net118));
 sg13g2_buf_8 fanout119 (.A(net121),
    .X(net119));
 sg13g2_buf_8 fanout120 (.A(net121),
    .X(net120));
 sg13g2_buf_8 fanout121 (.A(net122),
    .X(net121));
 sg13g2_buf_8 fanout122 (.A(_0824_),
    .X(net122));
 sg13g2_buf_8 fanout123 (.A(net124),
    .X(net123));
 sg13g2_buf_1 fanout124 (.A(_0823_),
    .X(net124));
 sg13g2_buf_8 fanout125 (.A(net127),
    .X(net125));
 sg13g2_buf_8 fanout126 (.A(net127),
    .X(net126));
 sg13g2_buf_8 fanout127 (.A(_0823_),
    .X(net127));
 sg13g2_buf_8 fanout128 (.A(net129),
    .X(net128));
 sg13g2_buf_8 fanout129 (.A(_0527_),
    .X(net129));
 sg13g2_buf_8 fanout130 (.A(_0482_),
    .X(net130));
 sg13g2_buf_8 fanout131 (.A(_0482_),
    .X(net131));
 sg13g2_buf_8 fanout132 (.A(_0437_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_0437_),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(_0392_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_0392_),
    .X(net135));
 sg13g2_buf_8 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_8 fanout137 (.A(_0347_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_1 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_8 fanout140 (.A(net141),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(net907),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(net143),
    .X(net142));
 sg13g2_buf_1 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(_0765_),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(_0765_),
    .X(net145));
 sg13g2_buf_8 fanout146 (.A(_0983_),
    .X(net146));
 sg13g2_buf_8 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(net898),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_1 fanout150 (.A(net900),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(net896),
    .X(net151));
 sg13g2_buf_8 fanout152 (.A(net892),
    .X(net152));
 sg13g2_buf_8 fanout153 (.A(net897),
    .X(net153));
 sg13g2_buf_8 fanout154 (.A(net899),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(net799),
    .X(net155));
 sg13g2_buf_8 fanout156 (.A(\u_cnt0.count[4] ),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(net160),
    .X(net157));
 sg13g2_buf_8 fanout158 (.A(net160),
    .X(net158));
 sg13g2_buf_8 fanout159 (.A(net160),
    .X(net159));
 sg13g2_buf_8 fanout160 (.A(_0960_),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(net167),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(net167),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(net167),
    .X(net164));
 sg13g2_buf_8 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_8 fanout167 (.A(rst_n),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(net173),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(net171),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(net173),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(rst_n),
    .X(net173));
 sg13g2_buf_1 input1 (.A(ui_in[2]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[3]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[4]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[5]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[6]),
    .X(net5));
 sg13g2_tielo tt_um_piggy_top_6 (.L_LO(net6));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_4 clkload4 (.A(clknet_leaf_42_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_leaf_43_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_0_clk));
 sg13g2_inv_2 clkload7 (.A(clknet_leaf_1_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_38_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_32_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_leaf_34_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_leaf_28_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_leaf_6_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_8_clk));
 sg13g2_inv_2 clkload14 (.A(clknet_leaf_9_clk));
 sg13g2_inv_2 clkload15 (.A(clknet_leaf_16_clk));
 sg13g2_inv_2 clkload16 (.A(clknet_leaf_22_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_25_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u_n2a2.ones[1] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold2 (.A(\u_n2a2.ones[0] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold3 (.A(\u_n2a0.ones[3] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold4 (.A(\u_n2a0.ones[0] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold5 (.A(\u_n2a3.ones[1] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold6 (.A(\u_n2a2.ones[3] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold7 (.A(\u_n2a2.ones[2] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold8 (.A(\u_n2a0.ones[1] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold9 (.A(\u_n2a3.ones[2] ),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u_n2a1.ones[0] ),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold11 (.A(\u_n2a3.ones[3] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u_n2a0.ones[2] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold13 (.A(\u_n2a1.ones[1] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold14 (.A(\u_n2a1.ones[3] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold15 (.A(\u_n2a1.ones[2] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold16 (.A(\u_n2a3.ones[0] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold17 (.A(\u_cnt3.count[0] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold18 (.A(\u_cnt2.count[0] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold19 (.A(\u_cnt1.count[0] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold20 (.A(\u_cnt0.count[0] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold21 (.A(\u_edge.state ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0154_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold23 (.A(\u_cnt1.state ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0123_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold25 (.A(\u_cnt2.state ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0133_),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u_cnt3.state ),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0143_),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold29 (.A(\u_cnt0.state ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0114_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold31 (.A(\u_n2a3.hundreds[0] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold32 (.A(\u_n2a2.hundreds[0] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u_n2a1.tens[1] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold34 (.A(\u_deb0.counter[0] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0009_),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold36 (.A(\u_n2a2.tens[2] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold37 (.A(\u_n2a1.tens[3] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold38 (.A(\u_deb4.counter[0] ),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0093_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold40 (.A(\u_n2a1.hundreds[0] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold41 (.A(\u_n2a3.hundreds[1] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold42 (.A(\u_n2a3.tens[3] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold43 (.A(\u_n2a1.tens[2] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold44 (.A(\u_n2a2.tens[3] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u_deb3.counter[0] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0072_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold47 (.A(\u_n2a2.tens[1] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold48 (.A(\u_n2a0.tens[2] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold49 (.A(\u_n2a0.hundreds[1] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold50 (.A(\u_n2a3.tens[2] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold51 (.A(\u_n2a0.tens[1] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold52 (.A(\u_deb1.counter[0] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0030_),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold54 (.A(\u_n2a0.hundreds[0] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold55 (.A(\u_n2a2.hundreds[1] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold56 (.A(\u_n2a1.hundreds[1] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold57 (.A(\u_n2a0.tens[3] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold58 (.A(\u_deb2.counter[0] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0051_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold60 (.A(\u_n2a2.tens[0] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold61 (.A(\u_n2a0.tens[0] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold62 (.A(\u_n2a3.tens[1] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold63 (.A(\u_uart.uart_tx_inst.clk_count[14] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold64 (.A(\u_uart.uart_tx_inst.clk_count[26] ),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold65 (.A(\u_uart.uart_tx_inst.clk_count[22] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0220_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold67 (.A(\u_uart.uart_tx_inst.clk_count[12] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold68 (.A(\u_uart.uart_tx_inst.clk_count[24] ),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0222_),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold70 (.A(\u_uart.uart_tx_inst.clk_count[27] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold71 (.A(\u_uart.uart_tx_inst.clk_count[19] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0217_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold73 (.A(\u_uart.uart_tx_inst.clk_count[20] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0218_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold75 (.A(\u_uart.uart_tx_inst.clk_count[11] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold76 (.A(\u_uart.uart_tx_inst.clk_count[16] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold77 (.A(\u_uart.uart_tx_inst.clk_count[25] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0223_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold79 (.A(\u_uart.uart_tx_inst.clk_count[31] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold80 (.A(\u_n2a3.tens[0] ),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold81 (.A(\u_uart.uart_tx_inst.clk_count[28] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold82 (.A(\u_uart.uart_tx_inst.clk_count[30] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold83 (.A(\u_uart.uart_tx_inst.clk_count[18] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0216_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold85 (.A(\u_n2a1.tens[0] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold86 (.A(\u_uart.uart_tx_inst.clk_count[17] ),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold87 (.A(\u_uart.uart_tx_inst.clk_count[23] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0221_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold89 (.A(\u_uart.uart_tx_inst.clk_count[21] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0219_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold91 (.A(\u_uart.uart_tx_inst.clk_count[15] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold92 (.A(\u_deb4.counter[18] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0559_),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0111_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold95 (.A(\u_uart.uart_tx_inst.clk_count[29] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold96 (.A(\u_deb4.counter[5] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0098_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold98 (.A(\u_deb0.counter[18] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0379_),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0027_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold101 (.A(\u_uart.uart_tx_inst.clk_count[13] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold102 (.A(\u_deb1.counter[5] ),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0035_),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold104 (.A(\u_deb2.counter[5] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0056_),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold106 (.A(\u_deb3.counter[18] ),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0514_),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0090_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold109 (.A(\u_deb0.counter[5] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0014_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold111 (.A(\u_deb3.counter[5] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0077_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold113 (.A(\u_deb1.counter[18] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0424_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0048_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold116 (.A(\u_deb2.counter[18] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0469_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0069_),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold119 (.A(\u_deb3.counter[6] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0492_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0078_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold122 (.A(\u_deb4.counter[6] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0537_),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0099_),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold125 (.A(\u_uart.uart_tx_inst.bit_index[2] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0232_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold127 (.A(\u_deb1.counter[6] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0402_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0036_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold130 (.A(\u_uart.uart_tx_inst.state[1] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0005_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold132 (.A(\u_deb0.counter[6] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0357_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0015_),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold135 (.A(\u_deb1.counter[17] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold136 (.A(_0047_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold137 (.A(\u_uart.state[3] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0235_),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold139 (.A(\u_deb3.counter[17] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0089_),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold141 (.A(\u_deb0.counter[17] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0026_),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold143 (.A(\u_deb4.counter[17] ),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0110_),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold145 (.A(\u_deb2.counter[17] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0068_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold147 (.A(\u_deb2.counter[6] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0447_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0057_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold150 (.A(\u_uart.uart_tx_inst.state[4] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold151 (.A(\u_uart.uart_tx_inst.clk_count[4] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0202_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold153 (.A(\u_uart.uart_tx_inst.clk_count[10] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0208_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold155 (.A(\u_uart.uart_tx_inst.tx_data[5] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0762_),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold157 (.A(\u_deb3.counter[2] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0485_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0074_),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold160 (.A(\u_cnt2.count[1] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0601_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold162 (.A(\u_deb2.Output ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold163 (.A(\u_deb2.counter[2] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0440_),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0053_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold166 (.A(\u_deb4.counter[2] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0530_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0095_),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold169 (.A(\u_deb1.counter[2] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0395_),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0032_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold172 (.A(\u_deb3.Output ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold173 (.A(\u_deb0.counter[2] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0350_),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0011_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold176 (.A(\u_cnt3.count[1] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold177 (.A(\u_deb4.Output ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold178 (.A(\u_deb0.Output ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold179 (.A(or4_out),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0635_),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold181 (.A(\u_uart.rom.addr[18] ),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0879_),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0254_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold184 (.A(\u_cnt1.count[1] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0283_),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold186 (.A(\u_uart.rom.addr[15] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0870_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0251_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold189 (.A(\u_deb2.counter[12] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0458_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0063_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold192 (.A(\u_deb0.counter[10] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0366_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0019_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold195 (.A(o_Tx_Done),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0000_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold197 (.A(\u_deb3.counter[12] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0503_),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0084_),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold200 (.A(\u_uart.rom.addr[13] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0249_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold202 (.A(\u_uart.rom.addr[12] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0860_),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0248_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold205 (.A(\u_deb1.counter[7] ),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0405_),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0037_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold208 (.A(\u_deb1.counter[3] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0398_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0033_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold211 (.A(\u_deb3.counter[3] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0488_),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0075_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold214 (.A(\u_deb4.counter[10] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0546_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0103_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold217 (.A(\u_deb1.counter[12] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0413_),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0042_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold220 (.A(\u_deb4.counter[3] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0533_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0096_),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold223 (.A(\u_deb0.counter[3] ),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0353_),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold225 (.A(_0012_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold226 (.A(\u_uart.rom.addr[9] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0850_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0245_),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold229 (.A(\u_uart.uart_tx_inst.clk_count[9] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0800_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0207_),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold232 (.A(\u_deb0.counter[12] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0368_),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0021_),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold235 (.A(\u_cnt0.count[1] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold236 (.A(\u_deb4.counter[12] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0548_),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0105_),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold239 (.A(\u_deb2.counter[7] ),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0450_),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0058_),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold242 (.A(\u_deb2.counter[3] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0443_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0054_),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold245 (.A(\u_deb0.counter[7] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0360_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold247 (.A(\u_deb2.counter[10] ),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0456_),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0061_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold250 (.A(\u_deb4.counter[7] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0540_),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold252 (.A(_0100_),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold253 (.A(\u_deb3.counter[9] ),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold254 (.A(_0498_),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0081_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold256 (.A(\u_deb4.counter[9] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0543_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0102_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold259 (.A(\u_deb4.counter[8] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0541_),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0101_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold262 (.A(\u_deb4.counter[4] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0534_),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0097_),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold265 (.A(\u_deb0.counter[16] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0376_),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0025_),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold268 (.A(\u_deb3.counter[7] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0495_),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0079_),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold271 (.A(\u_deb1.counter[10] ),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold272 (.A(_0411_),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0040_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold274 (.A(\u_deb4.counter[1] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0094_),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold276 (.A(\u_uart.rom.addr[16] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0252_),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold278 (.A(\u_deb2.counter[8] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0451_),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0059_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold281 (.A(\u_deb1.counter[8] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0406_),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0038_),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold284 (.A(\u_deb2.counter[19] ),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0435_),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold286 (.A(\u_deb1.counter[9] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0039_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold288 (.A(\u_deb3.counter[16] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0511_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold290 (.A(_0088_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold291 (.A(\u_deb0.counter[4] ),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold292 (.A(\u_deb4.counter[16] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0556_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0109_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold295 (.A(\u_deb3.counter[10] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0501_),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0082_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold298 (.A(\u_deb2.counter[9] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold299 (.A(\u_deb1.counter[4] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0034_),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold301 (.A(\u_deb1.counter[1] ),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0031_),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold303 (.A(\u_uart.state[2] ),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0987_),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0003_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold306 (.A(\u_uart.uart_tx_inst.clk_count[1] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold307 (.A(_0778_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0199_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold309 (.A(\u_deb3.counter[19] ),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0480_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold311 (.A(_0092_),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold312 (.A(\u_uart.uart_tx_inst.state[2] ),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold313 (.A(_0980_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold314 (.A(\u_deb0.counter[8] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold315 (.A(_0017_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold316 (.A(\u_deb2.counter[4] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold317 (.A(o_Tx_Active),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0809_),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0233_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold320 (.A(\u_deb2.counter[1] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold321 (.A(\u_deb0.counter[19] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold322 (.A(_0345_),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0029_),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold324 (.A(\u_uart.rom.addr[23] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0259_),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold326 (.A(\u_deb2.counter[16] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0466_),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0067_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold329 (.A(\u_deb3.counter[1] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold330 (.A(\u_deb3.counter[8] ),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold331 (.A(\u_deb0.counter[9] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold332 (.A(\u_deb0.counter[1] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold333 (.A(\u_uart.rom.addr[21] ),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0890_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold335 (.A(\u_deb4.counter[19] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0525_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold337 (.A(\u_uart.rom.addr[10] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0854_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold339 (.A(\u_uart.uart_tx_inst.tx_data[1] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0709_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0190_),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold342 (.A(\u_deb1.counter[16] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0421_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0046_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold345 (.A(\u_uart.rom.addr[6] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0840_),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold347 (.A(_0242_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold348 (.A(\u_uart.uart_tx_inst.clk_count[0] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold349 (.A(_0198_),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold350 (.A(\u_uart.rom.addr[20] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold351 (.A(\u_uart.rom.addr[25] ),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0905_),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold353 (.A(\u_deb3.counter[4] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold354 (.A(\u_deb1.Output ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold355 (.A(\u_uart.uart_tx_inst.tx_data[6] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold356 (.A(_0764_),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0195_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold358 (.A(\u_uart.rom.addr[30] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0921_),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0266_),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold361 (.A(\u_uart.rom.addr[28] ),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0916_),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold363 (.A(\u_uart.rom.addr[19] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0255_),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold365 (.A(\u_uart.uart_tx_inst.tx_data[0] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0691_),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0189_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold368 (.A(\u_uart.rom.addr[22] ),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold369 (.A(\u_uart.uart_tx_inst.clk_count[5] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0203_),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold371 (.A(\u_uart.rom.addr[29] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0265_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold373 (.A(\u_deb0.counter[11] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0020_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold375 (.A(\u_uart.rom.addr[26] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0262_),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold377 (.A(\u_deb1.counter[11] ),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0041_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold379 (.A(\u_uart.uart_tx_inst.tx_data[3] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0735_),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold381 (.A(_0192_),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold382 (.A(\u_uart.uart_tx_inst.tx_data[4] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0746_),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold384 (.A(\u_uart.uart_tx_inst.tx_data[2] ),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0191_),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold386 (.A(\u_deb4.counter[11] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold387 (.A(\u_deb2.counter[11] ),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold388 (.A(\u_cnt1.count[3] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0587_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0127_),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold391 (.A(start_sending),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold392 (.A(_0962_),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold393 (.A(\u_uart.uart_tx_inst.clk_count[2] ),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0200_),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold395 (.A(\u_deb1.counter[14] ),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0418_),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold397 (.A(_0044_),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold398 (.A(change0),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0770_),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold400 (.A(\u_deb3.counter[14] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0508_),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0086_),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold403 (.A(\u_deb0.counter[13] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold404 (.A(\u_uart.rom.addr[7] ),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold405 (.A(_0243_),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold406 (.A(\u_deb2.counter[13] ),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold407 (.A(\u_deb2.counter[14] ),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold408 (.A(\u_deb3.counter[11] ),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold409 (.A(\u_uart.rom.addr[24] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold410 (.A(\u_deb0.counter[15] ),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0375_),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0024_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold413 (.A(\u_uart.rom.addr[27] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold414 (.A(\u_uart.uart_tx_inst.state[0] ),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0819_),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold416 (.A(\u_deb4.counter[14] ),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold417 (.A(_0553_),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0107_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold419 (.A(\u_deb3.counter[15] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold420 (.A(\u_cnt0.count[4] ),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0571_),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold422 (.A(_0119_),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold423 (.A(\u_deb1.counter[15] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold424 (.A(\u_deb1.counter[13] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold425 (.A(\u_uart.rom.addr[1] ),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold426 (.A(_0237_),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold427 (.A(\u_deb2.counter[15] ),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold428 (.A(\u_deb1.counter[19] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold429 (.A(\u_deb4.counter[13] ),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold430 (.A(\u_deb4.counter[15] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold431 (.A(\u_uart.uart_tx_inst.clk_count[7] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold432 (.A(_0794_),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold433 (.A(\u_deb0.counter[14] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold434 (.A(\u_deb3.counter[13] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold435 (.A(\u_uart.state[1] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0004_),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold437 (.A(\u_cnt2.count[5] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0609_),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold439 (.A(\u_uart.uart_tx_inst.state[3] ),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold440 (.A(\u_uart.uart_tx_inst.i_Tx_Start [0]),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold441 (.A(\u_cnt2.count[2] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold442 (.A(\u_cnt1.count[6] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0593_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0130_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold445 (.A(\u_cnt0.count[2] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold446 (.A(\u_cnt1.count[2] ),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold447 (.A(\u_uart.rom.addr[17] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0253_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold449 (.A(\u_cnt1.count[5] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0591_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold451 (.A(\u_uart.uart_tx_inst.bit_index[1] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0978_),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold453 (.A(\u_uart.rom.addr[4] ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold454 (.A(\u_uart.uart_tx_inst.clk_count[8] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold455 (.A(_0796_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0206_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold457 (.A(\u_uart.rom.addr[11] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold458 (.A(\u_cnt0.count[5] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold459 (.A(\u_cnt3.count[5] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0627_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0149_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold462 (.A(\u_cnt0.count[6] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold463 (.A(\u_cnt0.count[3] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold464 (.A(\u_cnt3.count[2] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold465 (.A(\u_cnt2.count[6] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold466 (.A(\u_uart.rom.addr[8] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold467 (.A(\u_cnt1.count[7] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold468 (.A(\u_uart.rom.addr[31] ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold469 (.A(\u_cnt2.count[3] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold470 (.A(\u_uart.rom.addr[14] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold471 (.A(\u_cnt1.count[2] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold472 (.A(\u_uart.uart_tx_inst.clk_count[3] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold473 (.A(\u_uart.uart_tx_inst.bit_index[0] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold474 (.A(\u_cnt0.count[7] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold475 (.A(\u_cnt2.count[7] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold476 (.A(\u_cnt1.count[4] ),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold477 (.A(\u_cnt3.count[7] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold478 (.A(_0632_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold479 (.A(\u_uart.uart_tx_inst.clk_count[6] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold480 (.A(\u_uart.rom.addr[5] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold481 (.A(\u_cnt3.count[4] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold482 (.A(_0148_),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold483 (.A(\u_cnt3.count[2] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold484 (.A(\u_uart.rom.addr[0] ),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold485 (.A(\u_cnt3.count[6] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold486 (.A(\u_cnt3.count[3] ),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold487 (.A(\u_uart.rom.addr[3] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold488 (.A(\u_cnt2.count[4] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold489 (.A(\u_uart.rom.addr[2] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold490 (.A(\u_cnt1.count[5] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold491 (.A(\u_cnt3.count[5] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold492 (.A(\u_cnt0.count[6] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold493 (.A(\u_deb3.counter[4] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold494 (.A(\u_uart.rom.addr[5] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold495 (.A(\u_uart.uart_tx_inst.state[4] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold496 (.A(_0771_),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold497 (.A(\u_deb2.counter[1] ),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold498 (.A(\u_deb0.counter[1] ),
    .X(net909));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_fill_2 FILLER_0_175 ();
 sg13g2_fill_1 FILLER_0_177 ();
 sg13g2_decap_8 FILLER_0_192 ();
 sg13g2_decap_4 FILLER_0_199 ();
 sg13g2_decap_8 FILLER_0_208 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_decap_8 FILLER_0_222 ();
 sg13g2_decap_8 FILLER_0_229 ();
 sg13g2_decap_8 FILLER_0_236 ();
 sg13g2_decap_8 FILLER_0_243 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_decap_8 FILLER_0_257 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_313 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_334 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_4 FILLER_0_404 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_fill_1 FILLER_1_140 ();
 sg13g2_decap_4 FILLER_1_168 ();
 sg13g2_decap_4 FILLER_1_181 ();
 sg13g2_fill_1 FILLER_1_185 ();
 sg13g2_fill_1 FILLER_1_226 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_fill_1 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_237 ();
 sg13g2_decap_8 FILLER_2_244 ();
 sg13g2_decap_8 FILLER_2_251 ();
 sg13g2_decap_8 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_265 ();
 sg13g2_decap_8 FILLER_2_272 ();
 sg13g2_decap_8 FILLER_2_279 ();
 sg13g2_decap_8 FILLER_2_286 ();
 sg13g2_decap_8 FILLER_2_293 ();
 sg13g2_decap_8 FILLER_2_300 ();
 sg13g2_decap_8 FILLER_2_307 ();
 sg13g2_decap_8 FILLER_2_314 ();
 sg13g2_decap_8 FILLER_2_321 ();
 sg13g2_decap_8 FILLER_2_328 ();
 sg13g2_decap_8 FILLER_2_335 ();
 sg13g2_decap_8 FILLER_2_342 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_fill_1 FILLER_3_140 ();
 sg13g2_decap_4 FILLER_3_172 ();
 sg13g2_fill_1 FILLER_3_219 ();
 sg13g2_decap_8 FILLER_3_247 ();
 sg13g2_decap_8 FILLER_3_254 ();
 sg13g2_decap_8 FILLER_3_261 ();
 sg13g2_decap_8 FILLER_3_268 ();
 sg13g2_decap_8 FILLER_3_275 ();
 sg13g2_decap_8 FILLER_3_282 ();
 sg13g2_decap_8 FILLER_3_289 ();
 sg13g2_decap_8 FILLER_3_296 ();
 sg13g2_decap_8 FILLER_3_303 ();
 sg13g2_decap_8 FILLER_3_310 ();
 sg13g2_decap_8 FILLER_3_317 ();
 sg13g2_decap_8 FILLER_3_324 ();
 sg13g2_decap_8 FILLER_3_331 ();
 sg13g2_decap_8 FILLER_3_338 ();
 sg13g2_decap_8 FILLER_3_345 ();
 sg13g2_decap_8 FILLER_3_352 ();
 sg13g2_decap_8 FILLER_3_359 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_decap_8 FILLER_3_373 ();
 sg13g2_decap_8 FILLER_3_380 ();
 sg13g2_decap_8 FILLER_3_387 ();
 sg13g2_decap_8 FILLER_3_394 ();
 sg13g2_decap_8 FILLER_3_401 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_fill_2 FILLER_4_140 ();
 sg13g2_fill_1 FILLER_4_142 ();
 sg13g2_fill_2 FILLER_4_179 ();
 sg13g2_decap_4 FILLER_4_185 ();
 sg13g2_decap_4 FILLER_4_218 ();
 sg13g2_decap_8 FILLER_4_249 ();
 sg13g2_decap_8 FILLER_4_256 ();
 sg13g2_decap_8 FILLER_4_263 ();
 sg13g2_decap_8 FILLER_4_270 ();
 sg13g2_decap_8 FILLER_4_277 ();
 sg13g2_decap_8 FILLER_4_284 ();
 sg13g2_decap_8 FILLER_4_291 ();
 sg13g2_decap_8 FILLER_4_298 ();
 sg13g2_decap_8 FILLER_4_305 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_decap_8 FILLER_4_328 ();
 sg13g2_decap_8 FILLER_4_335 ();
 sg13g2_decap_8 FILLER_4_342 ();
 sg13g2_decap_8 FILLER_4_349 ();
 sg13g2_decap_8 FILLER_4_356 ();
 sg13g2_decap_8 FILLER_4_363 ();
 sg13g2_decap_8 FILLER_4_370 ();
 sg13g2_decap_8 FILLER_4_377 ();
 sg13g2_decap_8 FILLER_4_384 ();
 sg13g2_decap_8 FILLER_4_391 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_fill_1 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_fill_2 FILLER_5_194 ();
 sg13g2_fill_2 FILLER_5_206 ();
 sg13g2_fill_1 FILLER_5_208 ();
 sg13g2_fill_2 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_246 ();
 sg13g2_decap_8 FILLER_5_253 ();
 sg13g2_decap_8 FILLER_5_260 ();
 sg13g2_decap_8 FILLER_5_267 ();
 sg13g2_decap_8 FILLER_5_274 ();
 sg13g2_decap_8 FILLER_5_281 ();
 sg13g2_fill_2 FILLER_5_288 ();
 sg13g2_fill_1 FILLER_5_290 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_4 FILLER_6_140 ();
 sg13g2_fill_2 FILLER_6_144 ();
 sg13g2_fill_1 FILLER_6_173 ();
 sg13g2_decap_4 FILLER_6_187 ();
 sg13g2_decap_4 FILLER_6_219 ();
 sg13g2_fill_2 FILLER_6_223 ();
 sg13g2_decap_8 FILLER_6_229 ();
 sg13g2_fill_1 FILLER_6_236 ();
 sg13g2_decap_8 FILLER_6_264 ();
 sg13g2_decap_8 FILLER_6_271 ();
 sg13g2_decap_8 FILLER_6_278 ();
 sg13g2_fill_1 FILLER_6_317 ();
 sg13g2_decap_8 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_352 ();
 sg13g2_decap_8 FILLER_6_359 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_fill_1 FILLER_7_154 ();
 sg13g2_fill_2 FILLER_7_239 ();
 sg13g2_fill_1 FILLER_7_255 ();
 sg13g2_decap_8 FILLER_7_268 ();
 sg13g2_decap_8 FILLER_7_275 ();
 sg13g2_fill_2 FILLER_7_282 ();
 sg13g2_fill_1 FILLER_7_284 ();
 sg13g2_fill_2 FILLER_7_298 ();
 sg13g2_fill_1 FILLER_7_300 ();
 sg13g2_fill_2 FILLER_7_310 ();
 sg13g2_fill_1 FILLER_7_312 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_4 FILLER_8_147 ();
 sg13g2_decap_4 FILLER_8_155 ();
 sg13g2_fill_2 FILLER_8_159 ();
 sg13g2_fill_2 FILLER_8_197 ();
 sg13g2_fill_1 FILLER_8_199 ();
 sg13g2_decap_8 FILLER_8_278 ();
 sg13g2_decap_4 FILLER_8_285 ();
 sg13g2_fill_2 FILLER_8_289 ();
 sg13g2_decap_8 FILLER_8_360 ();
 sg13g2_decap_8 FILLER_8_367 ();
 sg13g2_decap_8 FILLER_8_374 ();
 sg13g2_decap_8 FILLER_8_381 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_161 ();
 sg13g2_fill_2 FILLER_9_187 ();
 sg13g2_fill_1 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_203 ();
 sg13g2_fill_1 FILLER_9_214 ();
 sg13g2_fill_2 FILLER_9_233 ();
 sg13g2_fill_1 FILLER_9_235 ();
 sg13g2_decap_8 FILLER_9_282 ();
 sg13g2_decap_8 FILLER_9_289 ();
 sg13g2_fill_2 FILLER_9_296 ();
 sg13g2_fill_2 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_355 ();
 sg13g2_decap_8 FILLER_9_362 ();
 sg13g2_decap_8 FILLER_9_369 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_4 FILLER_10_161 ();
 sg13g2_fill_2 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_171 ();
 sg13g2_fill_2 FILLER_10_178 ();
 sg13g2_fill_1 FILLER_10_239 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_fill_1 FILLER_10_289 ();
 sg13g2_fill_1 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_fill_2 FILLER_11_188 ();
 sg13g2_fill_1 FILLER_11_190 ();
 sg13g2_fill_2 FILLER_11_200 ();
 sg13g2_fill_1 FILLER_11_202 ();
 sg13g2_fill_2 FILLER_11_253 ();
 sg13g2_fill_2 FILLER_11_278 ();
 sg13g2_fill_1 FILLER_11_307 ();
 sg13g2_decap_8 FILLER_11_358 ();
 sg13g2_decap_8 FILLER_11_365 ();
 sg13g2_decap_8 FILLER_11_372 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_8 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_fill_1 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_106 ();
 sg13g2_decap_8 FILLER_12_113 ();
 sg13g2_decap_8 FILLER_12_120 ();
 sg13g2_decap_8 FILLER_12_127 ();
 sg13g2_decap_8 FILLER_12_134 ();
 sg13g2_decap_8 FILLER_12_141 ();
 sg13g2_decap_8 FILLER_12_148 ();
 sg13g2_decap_4 FILLER_12_155 ();
 sg13g2_fill_2 FILLER_12_159 ();
 sg13g2_fill_2 FILLER_12_188 ();
 sg13g2_fill_1 FILLER_12_190 ();
 sg13g2_decap_4 FILLER_12_222 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_decap_8 FILLER_12_275 ();
 sg13g2_fill_2 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_284 ();
 sg13g2_fill_2 FILLER_12_289 ();
 sg13g2_fill_1 FILLER_12_291 ();
 sg13g2_fill_2 FILLER_12_311 ();
 sg13g2_fill_1 FILLER_12_322 ();
 sg13g2_fill_1 FILLER_12_341 ();
 sg13g2_decap_8 FILLER_12_360 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_374 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_4 FILLER_13_56 ();
 sg13g2_fill_1 FILLER_13_60 ();
 sg13g2_fill_1 FILLER_13_66 ();
 sg13g2_decap_8 FILLER_13_71 ();
 sg13g2_fill_2 FILLER_13_78 ();
 sg13g2_fill_1 FILLER_13_80 ();
 sg13g2_decap_8 FILLER_13_114 ();
 sg13g2_decap_8 FILLER_13_121 ();
 sg13g2_decap_8 FILLER_13_128 ();
 sg13g2_decap_8 FILLER_13_135 ();
 sg13g2_decap_8 FILLER_13_142 ();
 sg13g2_decap_8 FILLER_13_149 ();
 sg13g2_fill_1 FILLER_13_156 ();
 sg13g2_fill_2 FILLER_13_214 ();
 sg13g2_fill_2 FILLER_13_234 ();
 sg13g2_fill_2 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_267 ();
 sg13g2_decap_8 FILLER_13_274 ();
 sg13g2_decap_4 FILLER_13_281 ();
 sg13g2_fill_2 FILLER_13_289 ();
 sg13g2_fill_2 FILLER_13_299 ();
 sg13g2_fill_2 FILLER_13_328 ();
 sg13g2_fill_1 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_49 ();
 sg13g2_fill_1 FILLER_14_89 ();
 sg13g2_fill_1 FILLER_14_136 ();
 sg13g2_decap_8 FILLER_14_150 ();
 sg13g2_decap_4 FILLER_14_157 ();
 sg13g2_fill_1 FILLER_14_161 ();
 sg13g2_fill_1 FILLER_14_166 ();
 sg13g2_decap_8 FILLER_14_192 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_215 ();
 sg13g2_fill_2 FILLER_14_285 ();
 sg13g2_fill_1 FILLER_14_314 ();
 sg13g2_fill_2 FILLER_14_328 ();
 sg13g2_fill_1 FILLER_14_330 ();
 sg13g2_fill_1 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_4 FILLER_15_42 ();
 sg13g2_fill_2 FILLER_15_46 ();
 sg13g2_decap_4 FILLER_15_76 ();
 sg13g2_fill_2 FILLER_15_124 ();
 sg13g2_fill_1 FILLER_15_126 ();
 sg13g2_decap_4 FILLER_15_163 ();
 sg13g2_fill_1 FILLER_15_167 ();
 sg13g2_fill_1 FILLER_15_181 ();
 sg13g2_fill_1 FILLER_15_243 ();
 sg13g2_fill_1 FILLER_15_294 ();
 sg13g2_fill_1 FILLER_15_304 ();
 sg13g2_decap_8 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_4 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_55 ();
 sg13g2_fill_1 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_226 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_4 FILLER_16_245 ();
 sg13g2_fill_1 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_332 ();
 sg13g2_fill_1 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_4 FILLER_17_63 ();
 sg13g2_decap_4 FILLER_17_98 ();
 sg13g2_fill_2 FILLER_17_102 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_4 FILLER_17_133 ();
 sg13g2_fill_1 FILLER_17_137 ();
 sg13g2_decap_8 FILLER_17_151 ();
 sg13g2_fill_2 FILLER_17_158 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_fill_2 FILLER_17_208 ();
 sg13g2_decap_4 FILLER_17_228 ();
 sg13g2_fill_1 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_241 ();
 sg13g2_decap_4 FILLER_17_247 ();
 sg13g2_decap_4 FILLER_17_272 ();
 sg13g2_fill_1 FILLER_17_276 ();
 sg13g2_decap_4 FILLER_17_286 ();
 sg13g2_fill_1 FILLER_17_298 ();
 sg13g2_fill_1 FILLER_17_304 ();
 sg13g2_fill_2 FILLER_17_309 ();
 sg13g2_fill_1 FILLER_17_321 ();
 sg13g2_fill_2 FILLER_17_327 ();
 sg13g2_fill_1 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_353 ();
 sg13g2_decap_8 FILLER_17_360 ();
 sg13g2_decap_8 FILLER_17_367 ();
 sg13g2_decap_8 FILLER_17_374 ();
 sg13g2_decap_8 FILLER_17_381 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_decap_8 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_4 FILLER_18_56 ();
 sg13g2_fill_1 FILLER_18_72 ();
 sg13g2_fill_2 FILLER_18_80 ();
 sg13g2_fill_1 FILLER_18_82 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_fill_1 FILLER_18_139 ();
 sg13g2_decap_8 FILLER_18_153 ();
 sg13g2_decap_4 FILLER_18_160 ();
 sg13g2_fill_2 FILLER_18_164 ();
 sg13g2_fill_1 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_212 ();
 sg13g2_decap_8 FILLER_18_219 ();
 sg13g2_fill_1 FILLER_18_226 ();
 sg13g2_fill_2 FILLER_18_256 ();
 sg13g2_fill_1 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_271 ();
 sg13g2_decap_8 FILLER_18_278 ();
 sg13g2_decap_8 FILLER_18_285 ();
 sg13g2_decap_8 FILLER_18_292 ();
 sg13g2_decap_4 FILLER_18_299 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_4 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_39 ();
 sg13g2_fill_1 FILLER_19_46 ();
 sg13g2_decap_4 FILLER_19_52 ();
 sg13g2_fill_1 FILLER_19_73 ();
 sg13g2_fill_1 FILLER_19_113 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_4 FILLER_19_175 ();
 sg13g2_fill_2 FILLER_19_179 ();
 sg13g2_fill_2 FILLER_19_188 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_208 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_fill_1 FILLER_19_216 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_fill_1 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_4 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_89 ();
 sg13g2_decap_4 FILLER_20_96 ();
 sg13g2_decap_4 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_125 ();
 sg13g2_decap_4 FILLER_20_132 ();
 sg13g2_fill_2 FILLER_20_136 ();
 sg13g2_decap_8 FILLER_20_169 ();
 sg13g2_decap_4 FILLER_20_190 ();
 sg13g2_fill_2 FILLER_20_338 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_37 ();
 sg13g2_decap_4 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_46 ();
 sg13g2_fill_1 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_86 ();
 sg13g2_decap_8 FILLER_21_93 ();
 sg13g2_decap_8 FILLER_21_100 ();
 sg13g2_decap_4 FILLER_21_107 ();
 sg13g2_fill_1 FILLER_21_111 ();
 sg13g2_fill_2 FILLER_21_139 ();
 sg13g2_fill_1 FILLER_21_141 ();
 sg13g2_decap_8 FILLER_21_155 ();
 sg13g2_fill_2 FILLER_21_162 ();
 sg13g2_fill_1 FILLER_21_164 ();
 sg13g2_decap_8 FILLER_21_234 ();
 sg13g2_fill_2 FILLER_21_241 ();
 sg13g2_decap_4 FILLER_21_275 ();
 sg13g2_fill_1 FILLER_21_279 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_fill_2 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_44 ();
 sg13g2_fill_1 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_68 ();
 sg13g2_decap_8 FILLER_22_75 ();
 sg13g2_decap_8 FILLER_22_82 ();
 sg13g2_decap_8 FILLER_22_89 ();
 sg13g2_decap_4 FILLER_22_96 ();
 sg13g2_fill_1 FILLER_22_100 ();
 sg13g2_decap_8 FILLER_22_106 ();
 sg13g2_decap_8 FILLER_22_113 ();
 sg13g2_decap_8 FILLER_22_120 ();
 sg13g2_decap_4 FILLER_22_127 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_fill_2 FILLER_22_168 ();
 sg13g2_fill_1 FILLER_22_170 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_211 ();
 sg13g2_decap_4 FILLER_22_216 ();
 sg13g2_fill_1 FILLER_22_220 ();
 sg13g2_decap_4 FILLER_22_227 ();
 sg13g2_decap_8 FILLER_22_244 ();
 sg13g2_fill_2 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_275 ();
 sg13g2_decap_8 FILLER_22_282 ();
 sg13g2_fill_1 FILLER_22_293 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_373 ();
 sg13g2_decap_8 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_44 ();
 sg13g2_decap_8 FILLER_23_64 ();
 sg13g2_decap_8 FILLER_23_71 ();
 sg13g2_fill_2 FILLER_23_85 ();
 sg13g2_fill_1 FILLER_23_87 ();
 sg13g2_fill_2 FILLER_23_96 ();
 sg13g2_fill_1 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_116 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_fill_2 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_170 ();
 sg13g2_decap_8 FILLER_23_177 ();
 sg13g2_decap_4 FILLER_23_188 ();
 sg13g2_fill_2 FILLER_23_192 ();
 sg13g2_decap_4 FILLER_23_208 ();
 sg13g2_fill_1 FILLER_23_212 ();
 sg13g2_fill_1 FILLER_23_216 ();
 sg13g2_decap_8 FILLER_23_254 ();
 sg13g2_fill_1 FILLER_23_261 ();
 sg13g2_decap_8 FILLER_23_290 ();
 sg13g2_fill_1 FILLER_23_297 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_352 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_55 ();
 sg13g2_fill_1 FILLER_24_57 ();
 sg13g2_decap_4 FILLER_24_75 ();
 sg13g2_fill_2 FILLER_24_90 ();
 sg13g2_fill_1 FILLER_24_111 ();
 sg13g2_fill_1 FILLER_24_139 ();
 sg13g2_decap_8 FILLER_24_153 ();
 sg13g2_decap_8 FILLER_24_160 ();
 sg13g2_fill_2 FILLER_24_167 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_decap_4 FILLER_24_230 ();
 sg13g2_fill_2 FILLER_24_261 ();
 sg13g2_fill_1 FILLER_24_263 ();
 sg13g2_decap_4 FILLER_24_273 ();
 sg13g2_fill_2 FILLER_24_277 ();
 sg13g2_fill_2 FILLER_24_284 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_fill_2 FILLER_24_368 ();
 sg13g2_fill_1 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_4 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_25 ();
 sg13g2_fill_2 FILLER_25_63 ();
 sg13g2_fill_1 FILLER_25_71 ();
 sg13g2_fill_1 FILLER_25_85 ();
 sg13g2_fill_1 FILLER_25_110 ();
 sg13g2_fill_1 FILLER_25_138 ();
 sg13g2_fill_1 FILLER_25_166 ();
 sg13g2_fill_1 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_25_234 ();
 sg13g2_decap_8 FILLER_25_257 ();
 sg13g2_fill_1 FILLER_25_264 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_42 ();
 sg13g2_fill_2 FILLER_26_46 ();
 sg13g2_fill_2 FILLER_26_74 ();
 sg13g2_fill_1 FILLER_26_76 ();
 sg13g2_decap_4 FILLER_26_111 ();
 sg13g2_fill_1 FILLER_26_115 ();
 sg13g2_fill_2 FILLER_26_170 ();
 sg13g2_fill_2 FILLER_26_279 ();
 sg13g2_fill_2 FILLER_26_300 ();
 sg13g2_fill_2 FILLER_26_338 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_33 ();
 sg13g2_fill_1 FILLER_27_35 ();
 sg13g2_fill_2 FILLER_27_55 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_69 ();
 sg13g2_fill_2 FILLER_27_85 ();
 sg13g2_fill_1 FILLER_27_87 ();
 sg13g2_decap_8 FILLER_27_100 ();
 sg13g2_decap_8 FILLER_27_107 ();
 sg13g2_decap_8 FILLER_27_118 ();
 sg13g2_fill_2 FILLER_27_125 ();
 sg13g2_fill_1 FILLER_27_132 ();
 sg13g2_fill_2 FILLER_27_146 ();
 sg13g2_fill_1 FILLER_27_148 ();
 sg13g2_decap_8 FILLER_27_157 ();
 sg13g2_decap_8 FILLER_27_164 ();
 sg13g2_decap_8 FILLER_27_171 ();
 sg13g2_decap_8 FILLER_27_178 ();
 sg13g2_fill_1 FILLER_27_185 ();
 sg13g2_decap_4 FILLER_27_191 ();
 sg13g2_decap_4 FILLER_27_204 ();
 sg13g2_fill_1 FILLER_27_208 ();
 sg13g2_decap_4 FILLER_27_213 ();
 sg13g2_fill_1 FILLER_27_217 ();
 sg13g2_fill_2 FILLER_27_305 ();
 sg13g2_fill_2 FILLER_27_311 ();
 sg13g2_fill_1 FILLER_27_313 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_21 ();
 sg13g2_fill_1 FILLER_28_23 ();
 sg13g2_fill_2 FILLER_28_52 ();
 sg13g2_fill_1 FILLER_28_54 ();
 sg13g2_decap_8 FILLER_28_90 ();
 sg13g2_decap_4 FILLER_28_97 ();
 sg13g2_decap_4 FILLER_28_104 ();
 sg13g2_fill_1 FILLER_28_108 ();
 sg13g2_decap_8 FILLER_28_136 ();
 sg13g2_decap_8 FILLER_28_170 ();
 sg13g2_decap_8 FILLER_28_177 ();
 sg13g2_decap_8 FILLER_28_184 ();
 sg13g2_decap_8 FILLER_28_191 ();
 sg13g2_decap_4 FILLER_28_198 ();
 sg13g2_fill_1 FILLER_28_202 ();
 sg13g2_decap_8 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_214 ();
 sg13g2_fill_2 FILLER_28_221 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_fill_2 FILLER_28_263 ();
 sg13g2_fill_2 FILLER_28_288 ();
 sg13g2_decap_8 FILLER_28_313 ();
 sg13g2_fill_2 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_322 ();
 sg13g2_decap_4 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_340 ();
 sg13g2_fill_1 FILLER_28_349 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_30 ();
 sg13g2_fill_2 FILLER_29_34 ();
 sg13g2_fill_1 FILLER_29_36 ();
 sg13g2_fill_1 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_75 ();
 sg13g2_fill_2 FILLER_29_82 ();
 sg13g2_decap_4 FILLER_29_87 ();
 sg13g2_fill_1 FILLER_29_91 ();
 sg13g2_decap_4 FILLER_29_128 ();
 sg13g2_decap_8 FILLER_29_145 ();
 sg13g2_decap_8 FILLER_29_152 ();
 sg13g2_decap_8 FILLER_29_159 ();
 sg13g2_fill_2 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_2 FILLER_29_254 ();
 sg13g2_fill_1 FILLER_29_256 ();
 sg13g2_decap_4 FILLER_29_261 ();
 sg13g2_fill_2 FILLER_29_276 ();
 sg13g2_fill_1 FILLER_29_295 ();
 sg13g2_fill_2 FILLER_29_310 ();
 sg13g2_fill_1 FILLER_29_312 ();
 sg13g2_decap_8 FILLER_29_335 ();
 sg13g2_decap_4 FILLER_29_342 ();
 sg13g2_fill_1 FILLER_29_346 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_4 FILLER_29_403 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_fill_2 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_30 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_4 FILLER_30_42 ();
 sg13g2_fill_1 FILLER_30_46 ();
 sg13g2_fill_1 FILLER_30_51 ();
 sg13g2_fill_1 FILLER_30_57 ();
 sg13g2_decap_8 FILLER_30_62 ();
 sg13g2_decap_4 FILLER_30_69 ();
 sg13g2_decap_8 FILLER_30_86 ();
 sg13g2_decap_4 FILLER_30_93 ();
 sg13g2_fill_2 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_167 ();
 sg13g2_fill_1 FILLER_30_196 ();
 sg13g2_fill_1 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_241 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_decap_4 FILLER_30_324 ();
 sg13g2_fill_1 FILLER_30_328 ();
 sg13g2_fill_2 FILLER_30_356 ();
 sg13g2_fill_2 FILLER_30_367 ();
 sg13g2_fill_1 FILLER_30_369 ();
 sg13g2_fill_1 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_45 ();
 sg13g2_decap_8 FILLER_31_52 ();
 sg13g2_decap_8 FILLER_31_59 ();
 sg13g2_decap_8 FILLER_31_66 ();
 sg13g2_decap_8 FILLER_31_73 ();
 sg13g2_decap_8 FILLER_31_80 ();
 sg13g2_decap_8 FILLER_31_87 ();
 sg13g2_fill_1 FILLER_31_94 ();
 sg13g2_fill_2 FILLER_31_129 ();
 sg13g2_fill_1 FILLER_31_158 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_201 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_fill_2 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_237 ();
 sg13g2_fill_2 FILLER_31_252 ();
 sg13g2_fill_1 FILLER_31_254 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_fill_1 FILLER_31_281 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_fill_2 FILLER_32_36 ();
 sg13g2_fill_1 FILLER_32_38 ();
 sg13g2_decap_8 FILLER_32_51 ();
 sg13g2_decap_8 FILLER_32_58 ();
 sg13g2_fill_2 FILLER_32_65 ();
 sg13g2_fill_1 FILLER_32_67 ();
 sg13g2_decap_8 FILLER_32_76 ();
 sg13g2_decap_8 FILLER_32_83 ();
 sg13g2_decap_8 FILLER_32_90 ();
 sg13g2_decap_8 FILLER_32_97 ();
 sg13g2_decap_8 FILLER_32_104 ();
 sg13g2_fill_2 FILLER_32_111 ();
 sg13g2_decap_4 FILLER_32_152 ();
 sg13g2_fill_2 FILLER_32_156 ();
 sg13g2_decap_4 FILLER_32_162 ();
 sg13g2_fill_2 FILLER_32_166 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_decap_4 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_254 ();
 sg13g2_decap_8 FILLER_32_261 ();
 sg13g2_fill_2 FILLER_32_268 ();
 sg13g2_fill_1 FILLER_32_270 ();
 sg13g2_fill_2 FILLER_32_284 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_fill_1 FILLER_32_304 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_fill_1 FILLER_33_19 ();
 sg13g2_fill_2 FILLER_33_64 ();
 sg13g2_decap_4 FILLER_33_86 ();
 sg13g2_fill_2 FILLER_33_117 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_decap_8 FILLER_33_170 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_fill_1 FILLER_33_187 ();
 sg13g2_decap_8 FILLER_33_202 ();
 sg13g2_decap_8 FILLER_33_209 ();
 sg13g2_fill_1 FILLER_33_222 ();
 sg13g2_fill_1 FILLER_33_227 ();
 sg13g2_fill_1 FILLER_33_237 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_fill_2 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_281 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_1 FILLER_33_294 ();
 sg13g2_fill_2 FILLER_33_309 ();
 sg13g2_fill_1 FILLER_33_352 ();
 sg13g2_fill_2 FILLER_33_367 ();
 sg13g2_fill_1 FILLER_33_369 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_69 ();
 sg13g2_fill_2 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_151 ();
 sg13g2_decap_4 FILLER_34_158 ();
 sg13g2_decap_4 FILLER_34_228 ();
 sg13g2_fill_1 FILLER_34_232 ();
 sg13g2_fill_1 FILLER_34_264 ();
 sg13g2_decap_4 FILLER_34_325 ();
 sg13g2_fill_2 FILLER_34_346 ();
 sg13g2_fill_1 FILLER_34_370 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_4 ();
 sg13g2_fill_2 FILLER_35_33 ();
 sg13g2_fill_2 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_79 ();
 sg13g2_fill_1 FILLER_35_151 ();
 sg13g2_fill_2 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_225 ();
 sg13g2_decap_4 FILLER_35_232 ();
 sg13g2_fill_1 FILLER_35_236 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_fill_2 FILLER_35_268 ();
 sg13g2_fill_1 FILLER_35_270 ();
 sg13g2_fill_1 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_325 ();
 sg13g2_fill_1 FILLER_35_327 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_23 ();
 sg13g2_fill_2 FILLER_36_40 ();
 sg13g2_decap_4 FILLER_36_50 ();
 sg13g2_fill_1 FILLER_36_54 ();
 sg13g2_decap_8 FILLER_36_59 ();
 sg13g2_decap_4 FILLER_36_66 ();
 sg13g2_fill_1 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_75 ();
 sg13g2_decap_8 FILLER_36_81 ();
 sg13g2_fill_1 FILLER_36_88 ();
 sg13g2_fill_1 FILLER_36_125 ();
 sg13g2_decap_8 FILLER_36_134 ();
 sg13g2_fill_1 FILLER_36_141 ();
 sg13g2_fill_1 FILLER_36_169 ();
 sg13g2_fill_2 FILLER_36_215 ();
 sg13g2_fill_1 FILLER_36_217 ();
 sg13g2_fill_2 FILLER_36_249 ();
 sg13g2_fill_2 FILLER_36_292 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_fill_1 FILLER_36_329 ();
 sg13g2_fill_2 FILLER_36_334 ();
 sg13g2_fill_1 FILLER_36_350 ();
 sg13g2_fill_2 FILLER_36_365 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_48 ();
 sg13g2_fill_1 FILLER_37_55 ();
 sg13g2_decap_8 FILLER_37_59 ();
 sg13g2_fill_1 FILLER_37_66 ();
 sg13g2_decap_8 FILLER_37_94 ();
 sg13g2_decap_8 FILLER_37_101 ();
 sg13g2_decap_8 FILLER_37_108 ();
 sg13g2_fill_1 FILLER_37_115 ();
 sg13g2_decap_8 FILLER_37_120 ();
 sg13g2_decap_8 FILLER_37_127 ();
 sg13g2_decap_8 FILLER_37_134 ();
 sg13g2_decap_4 FILLER_37_141 ();
 sg13g2_fill_2 FILLER_37_145 ();
 sg13g2_decap_8 FILLER_37_151 ();
 sg13g2_fill_1 FILLER_37_158 ();
 sg13g2_fill_1 FILLER_37_244 ();
 sg13g2_fill_2 FILLER_37_271 ();
 sg13g2_fill_2 FILLER_37_292 ();
 sg13g2_decap_8 FILLER_37_316 ();
 sg13g2_fill_2 FILLER_37_323 ();
 sg13g2_fill_2 FILLER_37_352 ();
 sg13g2_fill_1 FILLER_37_363 ();
 sg13g2_decap_8 FILLER_37_391 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_decap_4 FILLER_37_405 ();
 sg13g2_decap_4 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_4 ();
 sg13g2_decap_8 FILLER_38_39 ();
 sg13g2_decap_8 FILLER_38_46 ();
 sg13g2_decap_8 FILLER_38_115 ();
 sg13g2_decap_8 FILLER_38_127 ();
 sg13g2_decap_8 FILLER_38_134 ();
 sg13g2_fill_2 FILLER_38_141 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_267 ();
 sg13g2_fill_2 FILLER_38_274 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_4 FILLER_38_287 ();
 sg13g2_fill_1 FILLER_38_291 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_307 ();
 sg13g2_decap_8 FILLER_38_314 ();
 sg13g2_decap_8 FILLER_38_321 ();
 sg13g2_decap_8 FILLER_38_328 ();
 sg13g2_decap_8 FILLER_38_335 ();
 sg13g2_fill_2 FILLER_38_367 ();
 sg13g2_fill_1 FILLER_38_369 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_4 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_36 ();
 sg13g2_decap_8 FILLER_39_43 ();
 sg13g2_decap_8 FILLER_39_50 ();
 sg13g2_decap_8 FILLER_39_57 ();
 sg13g2_decap_8 FILLER_39_64 ();
 sg13g2_fill_1 FILLER_39_71 ();
 sg13g2_decap_8 FILLER_39_80 ();
 sg13g2_decap_4 FILLER_39_87 ();
 sg13g2_fill_1 FILLER_39_91 ();
 sg13g2_fill_2 FILLER_39_128 ();
 sg13g2_fill_1 FILLER_39_161 ();
 sg13g2_fill_2 FILLER_39_194 ();
 sg13g2_fill_1 FILLER_39_196 ();
 sg13g2_fill_2 FILLER_39_210 ();
 sg13g2_fill_1 FILLER_39_212 ();
 sg13g2_fill_2 FILLER_39_274 ();
 sg13g2_fill_1 FILLER_39_276 ();
 sg13g2_decap_8 FILLER_39_300 ();
 sg13g2_decap_4 FILLER_39_307 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_336 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_fill_2 FILLER_40_16 ();
 sg13g2_decap_4 FILLER_40_27 ();
 sg13g2_fill_1 FILLER_40_31 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_4 FILLER_40_70 ();
 sg13g2_fill_1 FILLER_40_74 ();
 sg13g2_decap_8 FILLER_40_79 ();
 sg13g2_decap_8 FILLER_40_86 ();
 sg13g2_fill_2 FILLER_40_93 ();
 sg13g2_fill_1 FILLER_40_126 ();
 sg13g2_decap_4 FILLER_40_172 ();
 sg13g2_fill_2 FILLER_40_181 ();
 sg13g2_fill_1 FILLER_40_183 ();
 sg13g2_fill_2 FILLER_40_197 ();
 sg13g2_decap_4 FILLER_40_208 ();
 sg13g2_fill_1 FILLER_40_212 ();
 sg13g2_fill_1 FILLER_40_283 ();
 sg13g2_decap_8 FILLER_40_356 ();
 sg13g2_fill_1 FILLER_40_363 ();
 sg13g2_fill_2 FILLER_40_368 ();
 sg13g2_fill_1 FILLER_40_370 ();
 sg13g2_fill_1 FILLER_40_384 ();
 sg13g2_fill_1 FILLER_40_389 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_fill_2 FILLER_40_406 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_29 ();
 sg13g2_fill_1 FILLER_41_42 ();
 sg13g2_fill_2 FILLER_41_50 ();
 sg13g2_fill_1 FILLER_41_69 ();
 sg13g2_fill_2 FILLER_41_97 ();
 sg13g2_fill_1 FILLER_41_99 ();
 sg13g2_fill_1 FILLER_41_113 ();
 sg13g2_decap_8 FILLER_41_145 ();
 sg13g2_fill_1 FILLER_41_152 ();
 sg13g2_fill_1 FILLER_41_163 ();
 sg13g2_decap_8 FILLER_41_170 ();
 sg13g2_decap_4 FILLER_41_177 ();
 sg13g2_decap_4 FILLER_41_192 ();
 sg13g2_fill_2 FILLER_41_231 ();
 sg13g2_fill_2 FILLER_41_238 ();
 sg13g2_fill_2 FILLER_41_247 ();
 sg13g2_fill_1 FILLER_41_249 ();
 sg13g2_fill_1 FILLER_41_305 ();
 sg13g2_decap_8 FILLER_41_338 ();
 sg13g2_decap_8 FILLER_41_345 ();
 sg13g2_fill_2 FILLER_41_366 ();
 sg13g2_fill_2 FILLER_41_392 ();
 sg13g2_fill_1 FILLER_41_394 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_12 ();
 sg13g2_fill_1 FILLER_42_14 ();
 sg13g2_fill_1 FILLER_42_41 ();
 sg13g2_decap_4 FILLER_42_68 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_127 ();
 sg13g2_decap_8 FILLER_42_134 ();
 sg13g2_decap_8 FILLER_42_141 ();
 sg13g2_decap_8 FILLER_42_148 ();
 sg13g2_decap_8 FILLER_42_155 ();
 sg13g2_decap_8 FILLER_42_167 ();
 sg13g2_fill_2 FILLER_42_174 ();
 sg13g2_fill_1 FILLER_42_176 ();
 sg13g2_fill_1 FILLER_42_199 ();
 sg13g2_fill_2 FILLER_42_240 ();
 sg13g2_fill_1 FILLER_42_242 ();
 sg13g2_fill_1 FILLER_42_292 ();
 sg13g2_fill_2 FILLER_42_298 ();
 sg13g2_fill_2 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_341 ();
 sg13g2_fill_1 FILLER_42_357 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_29 ();
 sg13g2_fill_2 FILLER_43_50 ();
 sg13g2_decap_8 FILLER_43_69 ();
 sg13g2_fill_1 FILLER_43_76 ();
 sg13g2_decap_8 FILLER_43_81 ();
 sg13g2_decap_8 FILLER_43_88 ();
 sg13g2_decap_8 FILLER_43_95 ();
 sg13g2_fill_2 FILLER_43_102 ();
 sg13g2_fill_1 FILLER_43_104 ();
 sg13g2_fill_2 FILLER_43_127 ();
 sg13g2_fill_2 FILLER_43_156 ();
 sg13g2_fill_1 FILLER_43_158 ();
 sg13g2_decap_4 FILLER_43_165 ();
 sg13g2_decap_8 FILLER_43_174 ();
 sg13g2_fill_1 FILLER_43_181 ();
 sg13g2_decap_8 FILLER_43_195 ();
 sg13g2_decap_8 FILLER_43_202 ();
 sg13g2_decap_4 FILLER_43_209 ();
 sg13g2_fill_2 FILLER_43_213 ();
 sg13g2_decap_4 FILLER_43_228 ();
 sg13g2_fill_2 FILLER_43_232 ();
 sg13g2_fill_2 FILLER_43_321 ();
 sg13g2_fill_1 FILLER_43_323 ();
 sg13g2_fill_2 FILLER_43_333 ();
 sg13g2_fill_1 FILLER_43_335 ();
 sg13g2_fill_1 FILLER_43_377 ();
 sg13g2_fill_1 FILLER_43_392 ();
 sg13g2_fill_2 FILLER_43_407 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_16 ();
 sg13g2_fill_2 FILLER_44_45 ();
 sg13g2_fill_2 FILLER_44_52 ();
 sg13g2_fill_2 FILLER_44_58 ();
 sg13g2_fill_2 FILLER_44_68 ();
 sg13g2_fill_2 FILLER_44_101 ();
 sg13g2_decap_4 FILLER_44_157 ();
 sg13g2_decap_8 FILLER_44_167 ();
 sg13g2_decap_8 FILLER_44_174 ();
 sg13g2_decap_4 FILLER_44_181 ();
 sg13g2_fill_2 FILLER_44_185 ();
 sg13g2_fill_1 FILLER_44_191 ();
 sg13g2_decap_8 FILLER_44_195 ();
 sg13g2_decap_8 FILLER_44_202 ();
 sg13g2_decap_8 FILLER_44_209 ();
 sg13g2_fill_1 FILLER_44_216 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_fill_1 FILLER_44_238 ();
 sg13g2_fill_2 FILLER_44_243 ();
 sg13g2_fill_1 FILLER_44_245 ();
 sg13g2_fill_1 FILLER_44_268 ();
 sg13g2_decap_4 FILLER_44_273 ();
 sg13g2_fill_2 FILLER_44_277 ();
 sg13g2_fill_2 FILLER_44_311 ();
 sg13g2_fill_1 FILLER_44_381 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_8 ();
 sg13g2_fill_1 FILLER_45_15 ();
 sg13g2_decap_4 FILLER_45_25 ();
 sg13g2_fill_1 FILLER_45_29 ();
 sg13g2_decap_4 FILLER_45_44 ();
 sg13g2_fill_2 FILLER_45_48 ();
 sg13g2_decap_8 FILLER_45_54 ();
 sg13g2_fill_2 FILLER_45_127 ();
 sg13g2_fill_1 FILLER_45_176 ();
 sg13g2_fill_2 FILLER_45_182 ();
 sg13g2_decap_4 FILLER_45_205 ();
 sg13g2_fill_2 FILLER_45_209 ();
 sg13g2_fill_2 FILLER_45_226 ();
 sg13g2_decap_8 FILLER_45_237 ();
 sg13g2_decap_8 FILLER_45_244 ();
 sg13g2_fill_2 FILLER_45_251 ();
 sg13g2_fill_1 FILLER_45_253 ();
 sg13g2_fill_1 FILLER_45_317 ();
 sg13g2_decap_4 FILLER_45_403 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_4 ();
 sg13g2_fill_1 FILLER_46_26 ();
 sg13g2_decap_4 FILLER_46_43 ();
 sg13g2_fill_1 FILLER_46_74 ();
 sg13g2_fill_2 FILLER_46_79 ();
 sg13g2_fill_1 FILLER_46_81 ();
 sg13g2_fill_2 FILLER_46_99 ();
 sg13g2_fill_2 FILLER_46_122 ();
 sg13g2_fill_1 FILLER_46_124 ();
 sg13g2_fill_2 FILLER_46_158 ();
 sg13g2_fill_1 FILLER_46_160 ();
 sg13g2_fill_2 FILLER_46_167 ();
 sg13g2_fill_1 FILLER_46_169 ();
 sg13g2_fill_2 FILLER_46_203 ();
 sg13g2_fill_1 FILLER_46_205 ();
 sg13g2_decap_8 FILLER_46_239 ();
 sg13g2_fill_2 FILLER_46_246 ();
 sg13g2_fill_1 FILLER_46_261 ();
 sg13g2_fill_2 FILLER_46_275 ();
 sg13g2_fill_1 FILLER_46_331 ();
 sg13g2_fill_1 FILLER_46_336 ();
 sg13g2_fill_1 FILLER_46_346 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_fill_2 FILLER_46_406 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_57 ();
 sg13g2_fill_1 FILLER_47_59 ();
 sg13g2_fill_1 FILLER_47_69 ();
 sg13g2_decap_8 FILLER_47_115 ();
 sg13g2_decap_8 FILLER_47_122 ();
 sg13g2_fill_1 FILLER_47_129 ();
 sg13g2_decap_8 FILLER_47_134 ();
 sg13g2_fill_2 FILLER_47_141 ();
 sg13g2_fill_1 FILLER_47_143 ();
 sg13g2_decap_8 FILLER_47_150 ();
 sg13g2_decap_8 FILLER_47_157 ();
 sg13g2_fill_2 FILLER_47_164 ();
 sg13g2_fill_1 FILLER_47_166 ();
 sg13g2_fill_1 FILLER_47_182 ();
 sg13g2_fill_1 FILLER_47_195 ();
 sg13g2_decap_4 FILLER_47_205 ();
 sg13g2_fill_2 FILLER_47_270 ();
 sg13g2_fill_2 FILLER_47_298 ();
 sg13g2_fill_2 FILLER_47_317 ();
 sg13g2_decap_4 FILLER_47_339 ();
 sg13g2_fill_2 FILLER_47_347 ();
 sg13g2_decap_8 FILLER_47_353 ();
 sg13g2_decap_4 FILLER_47_360 ();
 sg13g2_fill_2 FILLER_47_378 ();
 sg13g2_decap_4 FILLER_47_389 ();
 sg13g2_fill_1 FILLER_47_393 ();
 sg13g2_decap_4 FILLER_47_403 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_2 ();
 sg13g2_fill_2 FILLER_48_31 ();
 sg13g2_fill_1 FILLER_48_33 ();
 sg13g2_decap_8 FILLER_48_48 ();
 sg13g2_fill_2 FILLER_48_55 ();
 sg13g2_decap_8 FILLER_48_61 ();
 sg13g2_decap_8 FILLER_48_68 ();
 sg13g2_decap_8 FILLER_48_75 ();
 sg13g2_decap_8 FILLER_48_82 ();
 sg13g2_decap_8 FILLER_48_89 ();
 sg13g2_decap_8 FILLER_48_96 ();
 sg13g2_decap_8 FILLER_48_103 ();
 sg13g2_decap_4 FILLER_48_110 ();
 sg13g2_fill_1 FILLER_48_114 ();
 sg13g2_decap_8 FILLER_48_150 ();
 sg13g2_fill_2 FILLER_48_163 ();
 sg13g2_fill_1 FILLER_48_165 ();
 sg13g2_decap_8 FILLER_48_170 ();
 sg13g2_decap_4 FILLER_48_177 ();
 sg13g2_fill_2 FILLER_48_189 ();
 sg13g2_fill_1 FILLER_48_191 ();
 sg13g2_decap_8 FILLER_48_197 ();
 sg13g2_decap_8 FILLER_48_204 ();
 sg13g2_fill_2 FILLER_48_211 ();
 sg13g2_fill_2 FILLER_48_218 ();
 sg13g2_fill_2 FILLER_48_223 ();
 sg13g2_fill_1 FILLER_48_225 ();
 sg13g2_decap_4 FILLER_48_230 ();
 sg13g2_fill_1 FILLER_48_234 ();
 sg13g2_decap_8 FILLER_48_244 ();
 sg13g2_decap_8 FILLER_48_251 ();
 sg13g2_decap_8 FILLER_48_258 ();
 sg13g2_decap_4 FILLER_48_265 ();
 sg13g2_fill_2 FILLER_48_269 ();
 sg13g2_decap_8 FILLER_48_274 ();
 sg13g2_decap_4 FILLER_48_281 ();
 sg13g2_fill_1 FILLER_48_285 ();
 sg13g2_fill_2 FILLER_48_326 ();
 sg13g2_decap_8 FILLER_48_355 ();
 sg13g2_decap_8 FILLER_48_362 ();
 sg13g2_decap_8 FILLER_48_369 ();
 sg13g2_fill_1 FILLER_48_376 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_12 ();
 sg13g2_fill_2 FILLER_49_32 ();
 sg13g2_decap_8 FILLER_49_44 ();
 sg13g2_decap_8 FILLER_49_51 ();
 sg13g2_fill_1 FILLER_49_58 ();
 sg13g2_fill_2 FILLER_49_63 ();
 sg13g2_fill_1 FILLER_49_74 ();
 sg13g2_decap_4 FILLER_49_83 ();
 sg13g2_fill_2 FILLER_49_87 ();
 sg13g2_fill_2 FILLER_49_116 ();
 sg13g2_fill_2 FILLER_49_127 ();
 sg13g2_fill_2 FILLER_49_162 ();
 sg13g2_fill_1 FILLER_49_164 ();
 sg13g2_decap_4 FILLER_49_181 ();
 sg13g2_fill_2 FILLER_49_185 ();
 sg13g2_decap_8 FILLER_49_197 ();
 sg13g2_decap_8 FILLER_49_204 ();
 sg13g2_decap_8 FILLER_49_211 ();
 sg13g2_decap_8 FILLER_49_218 ();
 sg13g2_decap_8 FILLER_49_225 ();
 sg13g2_decap_8 FILLER_49_232 ();
 sg13g2_fill_1 FILLER_49_239 ();
 sg13g2_decap_4 FILLER_49_244 ();
 sg13g2_fill_2 FILLER_49_276 ();
 sg13g2_fill_1 FILLER_49_278 ();
 sg13g2_decap_8 FILLER_49_285 ();
 sg13g2_decap_4 FILLER_49_292 ();
 sg13g2_fill_2 FILLER_49_296 ();
 sg13g2_decap_4 FILLER_49_352 ();
 sg13g2_fill_2 FILLER_49_356 ();
 sg13g2_decap_8 FILLER_49_362 ();
 sg13g2_fill_2 FILLER_49_369 ();
 sg13g2_fill_1 FILLER_49_371 ();
 sg13g2_decap_4 FILLER_49_404 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_fill_1 FILLER_50_42 ();
 sg13g2_fill_2 FILLER_50_51 ();
 sg13g2_fill_1 FILLER_50_53 ();
 sg13g2_fill_2 FILLER_50_83 ();
 sg13g2_decap_4 FILLER_50_112 ();
 sg13g2_fill_1 FILLER_50_127 ();
 sg13g2_fill_2 FILLER_50_132 ();
 sg13g2_decap_8 FILLER_50_138 ();
 sg13g2_decap_8 FILLER_50_145 ();
 sg13g2_decap_4 FILLER_50_152 ();
 sg13g2_fill_2 FILLER_50_156 ();
 sg13g2_decap_8 FILLER_50_222 ();
 sg13g2_fill_2 FILLER_50_229 ();
 sg13g2_fill_2 FILLER_50_263 ();
 sg13g2_fill_1 FILLER_50_265 ();
 sg13g2_fill_1 FILLER_50_317 ();
 sg13g2_fill_2 FILLER_50_340 ();
 sg13g2_decap_8 FILLER_50_369 ();
 sg13g2_fill_1 FILLER_50_376 ();
 sg13g2_decap_4 FILLER_50_403 ();
 sg13g2_fill_2 FILLER_50_407 ();
 sg13g2_fill_1 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_29 ();
 sg13g2_fill_2 FILLER_51_49 ();
 sg13g2_fill_1 FILLER_51_51 ();
 sg13g2_fill_2 FILLER_51_60 ();
 sg13g2_fill_2 FILLER_51_72 ();
 sg13g2_fill_1 FILLER_51_74 ();
 sg13g2_decap_4 FILLER_51_80 ();
 sg13g2_fill_1 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_129 ();
 sg13g2_decap_8 FILLER_51_136 ();
 sg13g2_decap_8 FILLER_51_143 ();
 sg13g2_decap_8 FILLER_51_150 ();
 sg13g2_decap_8 FILLER_51_157 ();
 sg13g2_decap_8 FILLER_51_164 ();
 sg13g2_fill_2 FILLER_51_171 ();
 sg13g2_fill_1 FILLER_51_173 ();
 sg13g2_fill_2 FILLER_51_189 ();
 sg13g2_fill_1 FILLER_51_191 ();
 sg13g2_fill_1 FILLER_51_279 ();
 sg13g2_fill_1 FILLER_51_289 ();
 sg13g2_fill_1 FILLER_51_307 ();
 sg13g2_fill_2 FILLER_51_330 ();
 sg13g2_fill_1 FILLER_51_332 ();
 sg13g2_fill_2 FILLER_51_351 ();
 sg13g2_decap_4 FILLER_51_380 ();
 sg13g2_fill_1 FILLER_51_384 ();
 sg13g2_fill_2 FILLER_51_393 ();
 sg13g2_fill_1 FILLER_51_395 ();
 sg13g2_decap_4 FILLER_51_405 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_30 ();
 sg13g2_fill_2 FILLER_52_55 ();
 sg13g2_fill_1 FILLER_52_57 ();
 sg13g2_decap_8 FILLER_52_73 ();
 sg13g2_decap_8 FILLER_52_80 ();
 sg13g2_fill_2 FILLER_52_87 ();
 sg13g2_fill_1 FILLER_52_89 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_fill_2 FILLER_52_112 ();
 sg13g2_fill_2 FILLER_52_160 ();
 sg13g2_decap_8 FILLER_52_170 ();
 sg13g2_decap_4 FILLER_52_177 ();
 sg13g2_fill_2 FILLER_52_185 ();
 sg13g2_fill_1 FILLER_52_187 ();
 sg13g2_fill_1 FILLER_52_199 ();
 sg13g2_fill_2 FILLER_52_207 ();
 sg13g2_fill_1 FILLER_52_209 ();
 sg13g2_fill_2 FILLER_52_219 ();
 sg13g2_fill_1 FILLER_52_221 ();
 sg13g2_fill_1 FILLER_52_272 ();
 sg13g2_fill_2 FILLER_52_280 ();
 sg13g2_fill_1 FILLER_52_336 ();
 sg13g2_fill_1 FILLER_52_341 ();
 sg13g2_fill_2 FILLER_52_407 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_2 ();
 sg13g2_decap_4 FILLER_53_14 ();
 sg13g2_fill_1 FILLER_53_18 ();
 sg13g2_fill_2 FILLER_53_33 ();
 sg13g2_fill_2 FILLER_53_44 ();
 sg13g2_fill_1 FILLER_53_46 ();
 sg13g2_fill_1 FILLER_53_68 ();
 sg13g2_fill_2 FILLER_53_96 ();
 sg13g2_fill_2 FILLER_53_129 ();
 sg13g2_fill_1 FILLER_53_131 ();
 sg13g2_fill_2 FILLER_53_173 ();
 sg13g2_fill_1 FILLER_53_185 ();
 sg13g2_fill_1 FILLER_53_201 ();
 sg13g2_decap_8 FILLER_53_214 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_fill_1 FILLER_53_235 ();
 sg13g2_fill_1 FILLER_53_251 ();
 sg13g2_fill_1 FILLER_53_265 ();
 sg13g2_fill_2 FILLER_53_270 ();
 sg13g2_fill_2 FILLER_53_301 ();
 sg13g2_fill_1 FILLER_53_303 ();
 sg13g2_fill_2 FILLER_53_379 ();
 sg13g2_fill_1 FILLER_53_381 ();
 sg13g2_fill_2 FILLER_54_5 ();
 sg13g2_fill_1 FILLER_54_20 ();
 sg13g2_fill_1 FILLER_54_30 ();
 sg13g2_fill_1 FILLER_54_36 ();
 sg13g2_fill_2 FILLER_54_52 ();
 sg13g2_fill_1 FILLER_54_58 ();
 sg13g2_fill_1 FILLER_54_62 ();
 sg13g2_decap_4 FILLER_54_67 ();
 sg13g2_fill_2 FILLER_54_98 ();
 sg13g2_fill_1 FILLER_54_100 ();
 sg13g2_decap_8 FILLER_54_137 ();
 sg13g2_fill_1 FILLER_54_144 ();
 sg13g2_fill_2 FILLER_54_161 ();
 sg13g2_fill_1 FILLER_54_163 ();
 sg13g2_decap_4 FILLER_54_168 ();
 sg13g2_fill_2 FILLER_54_172 ();
 sg13g2_decap_4 FILLER_54_189 ();
 sg13g2_fill_1 FILLER_54_193 ();
 sg13g2_decap_8 FILLER_54_198 ();
 sg13g2_decap_4 FILLER_54_205 ();
 sg13g2_fill_1 FILLER_54_209 ();
 sg13g2_decap_8 FILLER_54_223 ();
 sg13g2_fill_1 FILLER_54_242 ();
 sg13g2_fill_1 FILLER_54_259 ();
 sg13g2_fill_1 FILLER_54_307 ();
 sg13g2_fill_2 FILLER_54_385 ();
 sg13g2_fill_2 FILLER_55_0 ();
 sg13g2_fill_2 FILLER_55_37 ();
 sg13g2_decap_8 FILLER_55_47 ();
 sg13g2_decap_8 FILLER_55_54 ();
 sg13g2_decap_8 FILLER_55_61 ();
 sg13g2_decap_4 FILLER_55_68 ();
 sg13g2_fill_1 FILLER_55_72 ();
 sg13g2_decap_8 FILLER_55_81 ();
 sg13g2_decap_8 FILLER_55_88 ();
 sg13g2_fill_1 FILLER_55_99 ();
 sg13g2_decap_8 FILLER_55_113 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_154 ();
 sg13g2_decap_8 FILLER_55_161 ();
 sg13g2_fill_2 FILLER_55_168 ();
 sg13g2_fill_1 FILLER_55_170 ();
 sg13g2_decap_4 FILLER_55_176 ();
 sg13g2_fill_2 FILLER_55_180 ();
 sg13g2_fill_1 FILLER_55_197 ();
 sg13g2_decap_8 FILLER_55_206 ();
 sg13g2_fill_2 FILLER_55_213 ();
 sg13g2_fill_2 FILLER_55_252 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_46 ();
 sg13g2_decap_4 FILLER_56_53 ();
 sg13g2_fill_2 FILLER_56_57 ();
 sg13g2_decap_8 FILLER_56_62 ();
 sg13g2_decap_8 FILLER_56_69 ();
 sg13g2_decap_8 FILLER_56_76 ();
 sg13g2_decap_4 FILLER_56_83 ();
 sg13g2_fill_2 FILLER_56_87 ();
 sg13g2_decap_8 FILLER_56_116 ();
 sg13g2_fill_2 FILLER_56_123 ();
 sg13g2_decap_8 FILLER_56_129 ();
 sg13g2_decap_8 FILLER_56_136 ();
 sg13g2_decap_8 FILLER_56_143 ();
 sg13g2_decap_8 FILLER_56_150 ();
 sg13g2_decap_8 FILLER_56_157 ();
 sg13g2_decap_8 FILLER_56_164 ();
 sg13g2_fill_1 FILLER_56_171 ();
 sg13g2_fill_2 FILLER_56_177 ();
 sg13g2_decap_8 FILLER_56_196 ();
 sg13g2_fill_1 FILLER_56_203 ();
 sg13g2_fill_1 FILLER_56_217 ();
 sg13g2_decap_8 FILLER_56_226 ();
 sg13g2_decap_4 FILLER_56_233 ();
 sg13g2_fill_2 FILLER_56_241 ();
 sg13g2_fill_1 FILLER_56_243 ();
 sg13g2_decap_8 FILLER_56_266 ();
 sg13g2_fill_2 FILLER_56_384 ();
 sg13g2_fill_1 FILLER_56_395 ();
 sg13g2_fill_1 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_50 ();
 sg13g2_decap_8 FILLER_57_57 ();
 sg13g2_fill_2 FILLER_57_64 ();
 sg13g2_decap_4 FILLER_57_71 ();
 sg13g2_decap_4 FILLER_57_91 ();
 sg13g2_fill_1 FILLER_57_95 ();
 sg13g2_decap_8 FILLER_57_100 ();
 sg13g2_fill_1 FILLER_57_134 ();
 sg13g2_decap_8 FILLER_57_181 ();
 sg13g2_decap_8 FILLER_57_188 ();
 sg13g2_decap_8 FILLER_57_195 ();
 sg13g2_fill_2 FILLER_57_202 ();
 sg13g2_decap_8 FILLER_57_218 ();
 sg13g2_fill_1 FILLER_57_241 ();
 sg13g2_decap_4 FILLER_57_259 ();
 sg13g2_fill_2 FILLER_57_272 ();
 sg13g2_fill_2 FILLER_57_291 ();
 sg13g2_fill_1 FILLER_57_298 ();
 sg13g2_fill_2 FILLER_57_334 ();
 sg13g2_fill_1 FILLER_57_336 ();
 sg13g2_fill_2 FILLER_57_383 ();
 sg13g2_fill_1 FILLER_57_385 ();
 sg13g2_decap_4 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_4 ();
 sg13g2_fill_1 FILLER_58_38 ();
 sg13g2_fill_2 FILLER_58_56 ();
 sg13g2_fill_2 FILLER_58_169 ();
 sg13g2_fill_1 FILLER_58_171 ();
 sg13g2_fill_2 FILLER_58_178 ();
 sg13g2_fill_1 FILLER_58_180 ();
 sg13g2_decap_8 FILLER_58_191 ();
 sg13g2_fill_1 FILLER_58_234 ();
 sg13g2_fill_2 FILLER_58_249 ();
 sg13g2_fill_1 FILLER_58_251 ();
 sg13g2_fill_2 FILLER_58_280 ();
 sg13g2_decap_8 FILLER_58_314 ();
 sg13g2_fill_2 FILLER_58_321 ();
 sg13g2_fill_1 FILLER_58_323 ();
 sg13g2_decap_8 FILLER_58_328 ();
 sg13g2_fill_2 FILLER_58_335 ();
 sg13g2_fill_1 FILLER_58_337 ();
 sg13g2_fill_2 FILLER_58_351 ();
 sg13g2_fill_1 FILLER_58_380 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_4 FILLER_59_19 ();
 sg13g2_fill_2 FILLER_59_45 ();
 sg13g2_fill_1 FILLER_59_47 ();
 sg13g2_decap_4 FILLER_59_88 ();
 sg13g2_decap_8 FILLER_59_96 ();
 sg13g2_fill_2 FILLER_59_147 ();
 sg13g2_fill_1 FILLER_59_149 ();
 sg13g2_decap_8 FILLER_59_163 ();
 sg13g2_decap_8 FILLER_59_170 ();
 sg13g2_decap_8 FILLER_59_177 ();
 sg13g2_fill_1 FILLER_59_215 ();
 sg13g2_decap_8 FILLER_59_278 ();
 sg13g2_fill_1 FILLER_59_285 ();
 sg13g2_fill_2 FILLER_59_299 ();
 sg13g2_fill_1 FILLER_59_301 ();
 sg13g2_decap_4 FILLER_59_311 ();
 sg13g2_fill_1 FILLER_59_360 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_20 ();
 sg13g2_fill_1 FILLER_60_29 ();
 sg13g2_fill_1 FILLER_60_54 ();
 sg13g2_decap_8 FILLER_60_76 ();
 sg13g2_decap_4 FILLER_60_83 ();
 sg13g2_fill_1 FILLER_60_114 ();
 sg13g2_decap_8 FILLER_60_137 ();
 sg13g2_fill_2 FILLER_60_144 ();
 sg13g2_fill_1 FILLER_60_146 ();
 sg13g2_decap_8 FILLER_60_182 ();
 sg13g2_decap_4 FILLER_60_193 ();
 sg13g2_fill_2 FILLER_60_197 ();
 sg13g2_fill_1 FILLER_60_226 ();
 sg13g2_fill_2 FILLER_60_236 ();
 sg13g2_fill_1 FILLER_60_238 ();
 sg13g2_fill_1 FILLER_60_266 ();
 sg13g2_decap_8 FILLER_60_280 ();
 sg13g2_decap_8 FILLER_60_287 ();
 sg13g2_decap_8 FILLER_60_294 ();
 sg13g2_decap_8 FILLER_60_301 ();
 sg13g2_decap_4 FILLER_60_308 ();
 sg13g2_fill_1 FILLER_60_312 ();
 sg13g2_fill_1 FILLER_60_318 ();
 sg13g2_fill_2 FILLER_60_324 ();
 sg13g2_fill_1 FILLER_60_326 ();
 sg13g2_fill_2 FILLER_60_381 ();
 sg13g2_fill_1 FILLER_60_383 ();
 sg13g2_fill_2 FILLER_60_398 ();
 sg13g2_decap_4 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_4 ();
 sg13g2_decap_4 FILLER_61_45 ();
 sg13g2_fill_2 FILLER_61_53 ();
 sg13g2_decap_8 FILLER_61_79 ();
 sg13g2_decap_8 FILLER_61_95 ();
 sg13g2_decap_8 FILLER_61_102 ();
 sg13g2_decap_8 FILLER_61_109 ();
 sg13g2_decap_4 FILLER_61_116 ();
 sg13g2_fill_2 FILLER_61_120 ();
 sg13g2_fill_2 FILLER_61_126 ();
 sg13g2_fill_1 FILLER_61_128 ();
 sg13g2_decap_8 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_185 ();
 sg13g2_decap_8 FILLER_61_192 ();
 sg13g2_fill_2 FILLER_61_199 ();
 sg13g2_decap_8 FILLER_61_218 ();
 sg13g2_fill_1 FILLER_61_225 ();
 sg13g2_decap_8 FILLER_61_230 ();
 sg13g2_fill_2 FILLER_61_237 ();
 sg13g2_decap_4 FILLER_61_246 ();
 sg13g2_fill_1 FILLER_61_250 ();
 sg13g2_fill_2 FILLER_61_256 ();
 sg13g2_fill_2 FILLER_61_271 ();
 sg13g2_fill_1 FILLER_61_273 ();
 sg13g2_decap_4 FILLER_61_278 ();
 sg13g2_fill_2 FILLER_61_282 ();
 sg13g2_fill_1 FILLER_61_311 ();
 sg13g2_fill_2 FILLER_61_384 ();
 sg13g2_fill_1 FILLER_61_386 ();
 sg13g2_fill_1 FILLER_61_396 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_fill_2 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_27 ();
 sg13g2_decap_8 FILLER_62_34 ();
 sg13g2_fill_2 FILLER_62_41 ();
 sg13g2_fill_1 FILLER_62_47 ();
 sg13g2_fill_2 FILLER_62_57 ();
 sg13g2_fill_1 FILLER_62_59 ();
 sg13g2_decap_8 FILLER_62_83 ();
 sg13g2_fill_2 FILLER_62_90 ();
 sg13g2_fill_1 FILLER_62_92 ();
 sg13g2_decap_8 FILLER_62_156 ();
 sg13g2_decap_8 FILLER_62_167 ();
 sg13g2_decap_8 FILLER_62_174 ();
 sg13g2_decap_8 FILLER_62_181 ();
 sg13g2_decap_8 FILLER_62_188 ();
 sg13g2_decap_8 FILLER_62_195 ();
 sg13g2_decap_8 FILLER_62_202 ();
 sg13g2_decap_8 FILLER_62_209 ();
 sg13g2_decap_8 FILLER_62_216 ();
 sg13g2_decap_4 FILLER_62_223 ();
 sg13g2_fill_1 FILLER_62_227 ();
 sg13g2_fill_1 FILLER_62_238 ();
 sg13g2_fill_2 FILLER_62_265 ();
 sg13g2_fill_1 FILLER_62_267 ();
 sg13g2_fill_1 FILLER_62_381 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_fill_2 FILLER_63_42 ();
 sg13g2_fill_1 FILLER_63_129 ();
 sg13g2_decap_8 FILLER_63_161 ();
 sg13g2_fill_1 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_209 ();
 sg13g2_decap_8 FILLER_63_216 ();
 sg13g2_fill_1 FILLER_63_223 ();
 sg13g2_decap_4 FILLER_63_269 ();
 sg13g2_fill_1 FILLER_63_273 ();
 sg13g2_fill_2 FILLER_63_288 ();
 sg13g2_fill_1 FILLER_63_290 ();
 sg13g2_fill_2 FILLER_63_313 ();
 sg13g2_fill_2 FILLER_63_377 ();
 sg13g2_fill_2 FILLER_63_389 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_fill_2 FILLER_64_21 ();
 sg13g2_fill_2 FILLER_64_86 ();
 sg13g2_fill_2 FILLER_64_115 ();
 sg13g2_fill_1 FILLER_64_117 ();
 sg13g2_fill_2 FILLER_64_136 ();
 sg13g2_fill_1 FILLER_64_138 ();
 sg13g2_decap_8 FILLER_64_143 ();
 sg13g2_fill_2 FILLER_64_150 ();
 sg13g2_fill_1 FILLER_64_152 ();
 sg13g2_fill_1 FILLER_64_180 ();
 sg13g2_decap_4 FILLER_64_221 ();
 sg13g2_fill_2 FILLER_64_318 ();
 sg13g2_fill_1 FILLER_64_320 ();
 sg13g2_fill_2 FILLER_64_398 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_fill_2 FILLER_65_21 ();
 sg13g2_fill_1 FILLER_65_23 ();
 sg13g2_fill_1 FILLER_65_33 ();
 sg13g2_fill_2 FILLER_65_62 ();
 sg13g2_fill_1 FILLER_65_64 ();
 sg13g2_decap_8 FILLER_65_74 ();
 sg13g2_fill_2 FILLER_65_81 ();
 sg13g2_fill_1 FILLER_65_83 ();
 sg13g2_decap_4 FILLER_65_96 ();
 sg13g2_fill_2 FILLER_65_100 ();
 sg13g2_fill_1 FILLER_65_106 ();
 sg13g2_decap_8 FILLER_65_111 ();
 sg13g2_decap_8 FILLER_65_118 ();
 sg13g2_decap_4 FILLER_65_125 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_4 FILLER_65_140 ();
 sg13g2_fill_1 FILLER_65_144 ();
 sg13g2_fill_1 FILLER_65_153 ();
 sg13g2_decap_4 FILLER_65_181 ();
 sg13g2_fill_1 FILLER_65_185 ();
 sg13g2_fill_1 FILLER_65_212 ();
 sg13g2_fill_2 FILLER_65_267 ();
 sg13g2_fill_1 FILLER_65_269 ();
 sg13g2_fill_2 FILLER_65_276 ();
 sg13g2_fill_1 FILLER_65_278 ();
 sg13g2_fill_1 FILLER_65_306 ();
 sg13g2_fill_2 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_fill_2 FILLER_66_28 ();
 sg13g2_fill_1 FILLER_66_30 ();
 sg13g2_decap_4 FILLER_66_48 ();
 sg13g2_decap_8 FILLER_66_61 ();
 sg13g2_fill_1 FILLER_66_68 ();
 sg13g2_decap_8 FILLER_66_73 ();
 sg13g2_decap_8 FILLER_66_80 ();
 sg13g2_decap_8 FILLER_66_87 ();
 sg13g2_decap_4 FILLER_66_94 ();
 sg13g2_fill_2 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_103 ();
 sg13g2_decap_8 FILLER_66_110 ();
 sg13g2_fill_2 FILLER_66_117 ();
 sg13g2_fill_1 FILLER_66_119 ();
 sg13g2_fill_1 FILLER_66_147 ();
 sg13g2_fill_2 FILLER_66_157 ();
 sg13g2_fill_1 FILLER_66_159 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_fill_1 FILLER_66_193 ();
 sg13g2_decap_8 FILLER_66_250 ();
 sg13g2_decap_4 FILLER_66_293 ();
 sg13g2_fill_2 FILLER_66_328 ();
 sg13g2_fill_1 FILLER_66_330 ();
 sg13g2_fill_1 FILLER_66_343 ();
 sg13g2_fill_2 FILLER_66_374 ();
 sg13g2_fill_1 FILLER_66_376 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_fill_2 FILLER_67_76 ();
 sg13g2_fill_1 FILLER_67_78 ();
 sg13g2_decap_8 FILLER_67_86 ();
 sg13g2_fill_1 FILLER_67_93 ();
 sg13g2_fill_2 FILLER_67_101 ();
 sg13g2_fill_1 FILLER_67_111 ();
 sg13g2_fill_2 FILLER_67_146 ();
 sg13g2_fill_1 FILLER_67_148 ();
 sg13g2_decap_4 FILLER_67_168 ();
 sg13g2_fill_1 FILLER_67_172 ();
 sg13g2_fill_2 FILLER_67_209 ();
 sg13g2_fill_1 FILLER_67_211 ();
 sg13g2_fill_1 FILLER_67_225 ();
 sg13g2_decap_4 FILLER_67_230 ();
 sg13g2_fill_1 FILLER_67_234 ();
 sg13g2_decap_8 FILLER_67_248 ();
 sg13g2_fill_2 FILLER_67_255 ();
 sg13g2_fill_1 FILLER_67_257 ();
 sg13g2_decap_8 FILLER_67_266 ();
 sg13g2_decap_8 FILLER_67_273 ();
 sg13g2_decap_4 FILLER_67_280 ();
 sg13g2_fill_1 FILLER_67_288 ();
 sg13g2_fill_2 FILLER_67_297 ();
 sg13g2_fill_1 FILLER_67_321 ();
 sg13g2_fill_2 FILLER_67_357 ();
 sg13g2_fill_1 FILLER_67_381 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_fill_2 FILLER_68_35 ();
 sg13g2_fill_1 FILLER_68_37 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_4 FILLER_68_49 ();
 sg13g2_fill_2 FILLER_68_53 ();
 sg13g2_fill_2 FILLER_68_70 ();
 sg13g2_fill_1 FILLER_68_72 ();
 sg13g2_fill_2 FILLER_68_114 ();
 sg13g2_fill_1 FILLER_68_116 ();
 sg13g2_decap_8 FILLER_68_134 ();
 sg13g2_fill_2 FILLER_68_141 ();
 sg13g2_fill_1 FILLER_68_143 ();
 sg13g2_decap_8 FILLER_68_175 ();
 sg13g2_fill_2 FILLER_68_182 ();
 sg13g2_decap_8 FILLER_68_220 ();
 sg13g2_decap_8 FILLER_68_227 ();
 sg13g2_fill_2 FILLER_68_234 ();
 sg13g2_fill_1 FILLER_68_236 ();
 sg13g2_decap_8 FILLER_68_242 ();
 sg13g2_decap_8 FILLER_68_249 ();
 sg13g2_fill_2 FILLER_68_256 ();
 sg13g2_decap_4 FILLER_68_271 ();
 sg13g2_fill_2 FILLER_68_275 ();
 sg13g2_fill_1 FILLER_68_304 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_fill_1 FILLER_69_32 ();
 sg13g2_fill_1 FILLER_69_61 ();
 sg13g2_fill_1 FILLER_69_81 ();
 sg13g2_fill_2 FILLER_69_87 ();
 sg13g2_fill_2 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_157 ();
 sg13g2_decap_8 FILLER_69_164 ();
 sg13g2_decap_8 FILLER_69_171 ();
 sg13g2_decap_8 FILLER_69_178 ();
 sg13g2_decap_4 FILLER_69_185 ();
 sg13g2_fill_2 FILLER_69_198 ();
 sg13g2_decap_8 FILLER_69_210 ();
 sg13g2_decap_8 FILLER_69_217 ();
 sg13g2_fill_1 FILLER_69_224 ();
 sg13g2_fill_1 FILLER_69_252 ();
 sg13g2_fill_2 FILLER_69_257 ();
 sg13g2_fill_1 FILLER_69_259 ();
 sg13g2_fill_1 FILLER_69_365 ();
 sg13g2_fill_2 FILLER_69_375 ();
 sg13g2_fill_1 FILLER_69_377 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_4 FILLER_70_14 ();
 sg13g2_fill_2 FILLER_70_18 ();
 sg13g2_fill_2 FILLER_70_51 ();
 sg13g2_decap_8 FILLER_70_90 ();
 sg13g2_fill_2 FILLER_70_97 ();
 sg13g2_decap_8 FILLER_70_104 ();
 sg13g2_decap_8 FILLER_70_115 ();
 sg13g2_decap_4 FILLER_70_122 ();
 sg13g2_decap_8 FILLER_70_130 ();
 sg13g2_decap_4 FILLER_70_137 ();
 sg13g2_fill_1 FILLER_70_141 ();
 sg13g2_fill_2 FILLER_70_209 ();
 sg13g2_fill_1 FILLER_70_265 ();
 sg13g2_fill_2 FILLER_70_270 ();
 sg13g2_fill_1 FILLER_70_282 ();
 sg13g2_fill_2 FILLER_70_302 ();
 sg13g2_fill_1 FILLER_70_330 ();
 sg13g2_fill_2 FILLER_70_354 ();
 sg13g2_fill_1 FILLER_70_383 ();
 sg13g2_fill_2 FILLER_70_397 ();
 sg13g2_fill_1 FILLER_70_399 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_fill_2 FILLER_71_21 ();
 sg13g2_fill_1 FILLER_71_23 ();
 sg13g2_fill_2 FILLER_71_53 ();
 sg13g2_fill_1 FILLER_71_55 ();
 sg13g2_fill_1 FILLER_71_65 ();
 sg13g2_fill_1 FILLER_71_70 ();
 sg13g2_fill_1 FILLER_71_75 ();
 sg13g2_fill_2 FILLER_71_114 ();
 sg13g2_decap_8 FILLER_71_120 ();
 sg13g2_fill_2 FILLER_71_127 ();
 sg13g2_fill_2 FILLER_71_172 ();
 sg13g2_fill_1 FILLER_71_230 ();
 sg13g2_fill_2 FILLER_71_249 ();
 sg13g2_fill_1 FILLER_71_251 ();
 sg13g2_fill_2 FILLER_71_274 ();
 sg13g2_fill_1 FILLER_71_276 ();
 sg13g2_fill_1 FILLER_71_309 ();
 sg13g2_fill_2 FILLER_71_328 ();
 sg13g2_fill_1 FILLER_71_330 ();
 sg13g2_fill_2 FILLER_71_345 ();
 sg13g2_fill_2 FILLER_71_370 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_fill_2 FILLER_72_40 ();
 sg13g2_fill_2 FILLER_72_47 ();
 sg13g2_fill_1 FILLER_72_49 ();
 sg13g2_fill_2 FILLER_72_54 ();
 sg13g2_fill_1 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_79 ();
 sg13g2_fill_2 FILLER_72_86 ();
 sg13g2_fill_2 FILLER_72_96 ();
 sg13g2_fill_2 FILLER_72_124 ();
 sg13g2_fill_2 FILLER_72_153 ();
 sg13g2_fill_1 FILLER_72_155 ();
 sg13g2_fill_1 FILLER_72_281 ();
 sg13g2_fill_2 FILLER_72_303 ();
 sg13g2_fill_1 FILLER_72_305 ();
 sg13g2_fill_1 FILLER_72_359 ();
 sg13g2_fill_2 FILLER_72_379 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_4 FILLER_73_21 ();
 sg13g2_fill_1 FILLER_73_25 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_fill_2 FILLER_73_121 ();
 sg13g2_fill_2 FILLER_73_131 ();
 sg13g2_fill_2 FILLER_73_277 ();
 sg13g2_fill_1 FILLER_73_279 ();
 sg13g2_fill_2 FILLER_73_321 ();
 sg13g2_fill_2 FILLER_73_350 ();
 sg13g2_fill_1 FILLER_73_352 ();
 sg13g2_fill_2 FILLER_73_367 ();
 sg13g2_fill_1 FILLER_73_369 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_fill_2 FILLER_74_28 ();
 sg13g2_fill_1 FILLER_74_30 ();
 sg13g2_decap_4 FILLER_74_35 ();
 sg13g2_fill_2 FILLER_74_76 ();
 sg13g2_fill_2 FILLER_74_83 ();
 sg13g2_decap_8 FILLER_74_94 ();
 sg13g2_decap_4 FILLER_74_101 ();
 sg13g2_fill_1 FILLER_74_105 ();
 sg13g2_fill_2 FILLER_74_127 ();
 sg13g2_decap_8 FILLER_74_173 ();
 sg13g2_decap_4 FILLER_74_180 ();
 sg13g2_fill_1 FILLER_74_184 ();
 sg13g2_fill_2 FILLER_74_198 ();
 sg13g2_fill_2 FILLER_74_213 ();
 sg13g2_fill_1 FILLER_74_215 ();
 sg13g2_fill_1 FILLER_74_221 ();
 sg13g2_fill_1 FILLER_74_259 ();
 sg13g2_fill_2 FILLER_74_304 ();
 sg13g2_fill_1 FILLER_74_306 ();
 sg13g2_fill_2 FILLER_74_316 ();
 sg13g2_fill_1 FILLER_74_323 ();
 sg13g2_fill_1 FILLER_74_345 ();
 sg13g2_fill_1 FILLER_74_382 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_4 FILLER_75_28 ();
 sg13g2_fill_2 FILLER_75_71 ();
 sg13g2_fill_1 FILLER_75_73 ();
 sg13g2_fill_1 FILLER_75_100 ();
 sg13g2_decap_8 FILLER_75_106 ();
 sg13g2_decap_8 FILLER_75_129 ();
 sg13g2_fill_2 FILLER_75_136 ();
 sg13g2_decap_4 FILLER_75_142 ();
 sg13g2_fill_1 FILLER_75_200 ();
 sg13g2_fill_2 FILLER_75_271 ();
 sg13g2_fill_1 FILLER_75_273 ();
 sg13g2_fill_1 FILLER_75_309 ();
 sg13g2_fill_2 FILLER_75_315 ();
 sg13g2_fill_1 FILLER_75_317 ();
 sg13g2_fill_2 FILLER_75_335 ();
 sg13g2_fill_2 FILLER_75_380 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_4 FILLER_76_21 ();
 sg13g2_fill_1 FILLER_76_25 ();
 sg13g2_fill_2 FILLER_76_44 ();
 sg13g2_fill_2 FILLER_76_55 ();
 sg13g2_fill_2 FILLER_76_62 ();
 sg13g2_fill_2 FILLER_76_69 ();
 sg13g2_fill_1 FILLER_76_71 ();
 sg13g2_decap_4 FILLER_76_82 ();
 sg13g2_fill_1 FILLER_76_86 ();
 sg13g2_decap_8 FILLER_76_96 ();
 sg13g2_decap_8 FILLER_76_103 ();
 sg13g2_decap_4 FILLER_76_110 ();
 sg13g2_decap_8 FILLER_76_122 ();
 sg13g2_decap_4 FILLER_76_129 ();
 sg13g2_fill_1 FILLER_76_133 ();
 sg13g2_decap_4 FILLER_76_138 ();
 sg13g2_fill_2 FILLER_76_142 ();
 sg13g2_fill_2 FILLER_76_157 ();
 sg13g2_decap_8 FILLER_76_163 ();
 sg13g2_decap_8 FILLER_76_170 ();
 sg13g2_fill_1 FILLER_76_177 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_fill_2 FILLER_76_189 ();
 sg13g2_fill_2 FILLER_76_237 ();
 sg13g2_fill_1 FILLER_76_239 ();
 sg13g2_fill_2 FILLER_76_281 ();
 sg13g2_fill_2 FILLER_76_348 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_65 ();
 sg13g2_fill_1 FILLER_77_72 ();
 sg13g2_decap_8 FILLER_77_82 ();
 sg13g2_fill_1 FILLER_77_89 ();
 sg13g2_fill_1 FILLER_77_100 ();
 sg13g2_decap_8 FILLER_77_106 ();
 sg13g2_fill_1 FILLER_77_113 ();
 sg13g2_fill_2 FILLER_77_123 ();
 sg13g2_fill_1 FILLER_77_125 ();
 sg13g2_fill_1 FILLER_77_153 ();
 sg13g2_decap_4 FILLER_77_181 ();
 sg13g2_fill_1 FILLER_77_185 ();
 sg13g2_fill_1 FILLER_77_297 ();
 sg13g2_fill_1 FILLER_77_361 ();
 sg13g2_fill_2 FILLER_77_384 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_4 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_76 ();
 sg13g2_fill_1 FILLER_78_83 ();
 sg13g2_decap_4 FILLER_78_127 ();
 sg13g2_decap_8 FILLER_78_135 ();
 sg13g2_fill_2 FILLER_78_142 ();
 sg13g2_fill_1 FILLER_78_144 ();
 sg13g2_decap_4 FILLER_78_149 ();
 sg13g2_fill_1 FILLER_78_153 ();
 sg13g2_decap_8 FILLER_78_163 ();
 sg13g2_decap_8 FILLER_78_170 ();
 sg13g2_fill_2 FILLER_78_177 ();
 sg13g2_fill_1 FILLER_78_225 ();
 sg13g2_fill_1 FILLER_78_239 ();
 sg13g2_fill_2 FILLER_78_346 ();
 sg13g2_fill_1 FILLER_78_381 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_4 FILLER_79_35 ();
 sg13g2_fill_1 FILLER_79_39 ();
 sg13g2_fill_2 FILLER_79_49 ();
 sg13g2_fill_1 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_167 ();
 sg13g2_decap_8 FILLER_79_174 ();
 sg13g2_decap_4 FILLER_79_181 ();
 sg13g2_fill_1 FILLER_79_185 ();
 sg13g2_fill_2 FILLER_79_270 ();
 sg13g2_fill_1 FILLER_79_317 ();
 sg13g2_fill_1 FILLER_79_380 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_fill_2 FILLER_80_49 ();
 sg13g2_fill_1 FILLER_80_51 ();
 sg13g2_fill_2 FILLER_80_60 ();
 sg13g2_fill_2 FILLER_80_70 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_fill_2 FILLER_80_125 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_fill_2 FILLER_80_149 ();
 sg13g2_fill_1 FILLER_80_151 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_4 FILLER_80_180 ();
 sg13g2_fill_1 FILLER_80_188 ();
 sg13g2_fill_2 FILLER_80_197 ();
 sg13g2_fill_1 FILLER_80_199 ();
 sg13g2_fill_2 FILLER_80_212 ();
 sg13g2_fill_1 FILLER_80_231 ();
 sg13g2_fill_1 FILLER_80_241 ();
 sg13g2_fill_2 FILLER_80_251 ();
 sg13g2_fill_2 FILLER_80_258 ();
 sg13g2_fill_1 FILLER_80_260 ();
 sg13g2_fill_2 FILLER_80_287 ();
 sg13g2_fill_1 FILLER_80_289 ();
 sg13g2_fill_1 FILLER_80_326 ();
 sg13g2_fill_2 FILLER_80_353 ();
 sg13g2_fill_1 FILLER_80_355 ();
 sg13g2_fill_1 FILLER_80_397 ();
 sg13g2_fill_2 FILLER_80_407 ();
 assign uio_oe[0] = net6;
 assign uio_oe[1] = net7;
 assign uio_oe[2] = net8;
 assign uio_oe[3] = net9;
 assign uio_oe[4] = net10;
 assign uio_oe[5] = net11;
 assign uio_oe[6] = net12;
 assign uio_oe[7] = net13;
 assign uio_out[0] = net14;
 assign uio_out[1] = net15;
 assign uio_out[2] = net16;
 assign uio_out[3] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
 assign uo_out[3] = net22;
 assign uo_out[4] = net23;
 assign uo_out[5] = net24;
 assign uo_out[6] = net25;
 assign uo_out[7] = net26;
endmodule
